��J     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.3.0�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh&hNhJ�
hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��h4�f8�����R�(KhQNNNJ����J����K t�b�C              �?�t�bhUh(�scalar���hPC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hK�
node_count�KՌnodes�h*h-K ��h/��R�(KKՅ�h4�V64�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h�hPK ��h�hPK��h�hPK��h�haK��h�haK ��h�hPK(��h�haK0��h�h4�u1�����R�(Kh8NNNJ����J����K t�bK8��uK@KKt�b�B@5         P                    �?j8je3�?�           ��@                                   �?���̟�?�            r@ A,160,3       
       
             �?X�If%��?\            �b@ \ u t                            �?�Ru߬Α?G            �\@ i g   ������������������������       �        @            @Y@               	                    @K@$�q-�?             *@                                  @d@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?
    >>>������������������������       �                     @fit([[-1              	             �?�t����?             A@ nonzero                           �?�z�G��?             $@  �bool������������������������       �                      @ndom_sta                           �?      �?              @o_coefs                           �D@z�G�z�?             @ r   FT������������������������       �                     �? _|| _������������������������       �                     @t,1
54,������������������������       �                     @                                   @L@      �?             8@                                   �?�z�G��?             $@B��fn                          �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @��`3���������������������������       �                     ,@               )                   �]@��t�?_            �a@               &                   �c@������?             ;@              %                   p`@�㙢�c�?             7@                                  �?����X�?
             ,@        ������������������������       �                     @                       	          fff�?���Q��?             $@        ������������������������       �                     @        !       "                   �c@؇���X�?             @ c t o ������������������������       �                     @M��b��#       $                    �?      �?              @        ������������������������       �                     �?D�:5ݠ�������������������������       �                     �?      _ ������������������������       �                     "@ex=['cat'       (       	             �?      �?             @   colum������������������������       �                     �?es when ������������������������       �                     @s the st*       I       	          pff�?���;�?N            �\@e origi+       @                    �?��!���?C            @W@s:

   ,       3       
             �?���?:            �R@       -       2                    �?@3����?(             K@  3.0  .       /                   �s@P�Lt�<�?             C@      h������������������������       �                     B@ m      0       1                    �N@      �?              @      4.������������������������       �                     �?ked**

 ������������������������       �                     �?s are st������������������������       �                     0@        4       9                    @K@�G��l��?             5@ eight  5       6                    ]@z�G�z�?             $@  3.0  N������������������������       �                     �?  cat  h7       8                   �q@�����H�?             "@og  hei������������������������       �                      @ype: flo������������������������       �                     �?f_multi_:       ;                   �p@���!pc�?
             &@     ..������������������������       �                     @'],
    <       ?                   �`@      �?             @col2)

=       >                    �?      �?              @ ropped ������������������������       �                     �?via the ������������������������       �                     �?level_co������������������������       �                      @        A       B                    l@X�<ݚ�?	             2@        ������������������������       �                      @      �?C       H                   �q@z�G�z�?             $@       D       E                    @M@�����H�?             "@       ������������������������       �                     @        F       G                    �P@      �?              @      �?������������������������       �                     �?      �?������������������������       �                     �?        ������������������������       �                     �?        J       O                   ``@���N8�?             5@     �?K       L                     G@�eP*L��?             &@        ������������������������       �                     @        M       N                   @_@      �?              @        ������������������������       �                     @      �?������������������������       �                      @      �?������������������������       �                     $@        Q       �                   a@�����L�?           �{@     �?R       c       
             �?�u2�dD�?�            �p@        S       Z                    �?      �?             @@        T       Y                    �?      �?             0@       U       V       	          hff�?z�G�z�?             $@       ������������������������       �                     @        W       X                    �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @      �?[       ^                   �W@      �?             0@      �?\       ]       	          @33�?      �?             @p�#�������������������������       �                     @�       ������������������������       �                     �?Z      _       b                    �E@�8��8��?
             (@       `       a                   �\@      �?              @       ������������������������       �                     �?N      ������������������������       �                     �?�       ������������������������       �                     $@�       d       e       	             �?l{��b��?�            �m@       ������������������������       �                    �I@�       f       g                   �Q@��a�n`�?v            @g@       ������������������������       �                      @      h       �                    @���}<S�?u             g@      i       �                    �?4����Y�?q            �e@      j       y                   `_@     �?U             `@      k       x                    �L@ p�/��?>            @V@      l       w                   �[@l�b�G��?&            �L@       m       v                   �a@PN��T'�?             ;@       n       u                    �?���|���?	             &@      o       t                    �?      �?              @      p       s                   �Z@և���X�?             @      q       r                    �K@      �?             @      ������������������������       �                     @�       ������������������������       �                     �?�      ������������������������       �                     @�      ������������������������       �                     �?�      ������������������������       �                     @P       ������������������������       �        
             0@�      ������������������������       �                     >@�      ������������������������       �                     @@       z       �                   p`@:�&���?            �C@       {       �       	          ����?R�}e�.�?             :@       |       }                   p`@�z�G��?             $@       ������������������������       �                     @�      ~                           l@      �?             @      ������������������������       �                     @�       ������������������������       �                     �?~      ������������������������       �        
             0@�       ������������������������       �                     *@�      �       �       
             �?`Ql�R�?            �G@       ������������������������       �                     C@g       �       �                   �[@�����H�?             "@       ������������������������       �                     @      �       �                   `c@z�G�z�?             @      ������������������������       �                     @�      ������������������������       �                     �?�      �       �                   �k@X�<ݚ�?             "@       ������������������������       �                     @�      ������������������������       �                     @�      �       �                   Pq@      �?l             f@      �       �       
             �?�ȋ}��?T            @`@       �       �                    �?^(��I�?&            �K@      �       �                    �?H.�!���?"             I@      �       �                    �?�(�Tw��?            �C@       �       �                   @e@�q�q�?             "@      ������������������������       �                     @      ������������������������       �                     @m      �       �                   pe@������?             >@       ������������������������       �                     @R      �       �                   �e@�q�q�?             8@       ������������������������       �                     �?�       �       �                   �p@8����?             7@       �       �                    �?��Q��?             4@       �       �                   �o@�n_Y�K�?
             *@       �       �                   l@���!pc�?	             &@       �       �                    @      �?             @       �       �                    j@���Q��?             @        ������������������������       �                      @�       �       �       	             �?�q�q�?             @       �       �                   �e@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?-       ������������������������       �                     �?_       ������������������������       �                     �?T       ������������������������       �                     @B       ������������������������       �                      @3       �       �                   �n@����X�?             @      ������������������������       �                     @�      ������������������������       �                      @w      ������������������������       �                     @j      ������������������������       �                     &@�      �       �                    �?���Q��?             @      ������������������������       �                     @�      ������������������������       �                      @�      �       �                   �Z@DE��2{�?.            �R@       �       �                    �?���Q��?             @      ������������������������       �                     @       ������������������������       �                      @�       �       �                    �?z��R[�?+            �Q@      �       �                    q@lGts��?"            �K@      �       �       	          033�?�NW���?!            �J@      �       �                    �?�J�4�?             9@      �       �       	          ����?����X�?             ,@ps �������������������������       �                     "@        �       �                   �g@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     <@        ������������������������       �                      @        �       �       	          ���@��S���?	             .@       �       �                    �?�<ݚ�?             "@        �       �                    _@      �?             @       �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     J@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @F@�3Ea�$�?             G@        �       �                   @_@      �?             ,@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �L@      �?             @@        �       �                    @L@؇���X�?             ,@       ������������������������       �                     &@        �       �       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             2@        �t�b�values�h*h-K ��h/��R�(KK�KK��ha�BP       Ps@     �z@      j@      T@     �^@      9@     @\@      �?     @Y@              (@      �?      @      �?      @                      �?      @              $@      8@      @      @               @      @      �?      @      �?              �?      @              @              @      5@      @      @      �?      @      �?                      @       @                      ,@     �U@     �K@      @      4@      @      3@      @      $@              @      @      @      @              �?      @              @      �?      �?              �?      �?                      "@      @      �?              �?      @             �S@     �A@     �R@      3@      P@      &@     �J@      �?     �B@      �?      B@              �?      �?      �?                      �?      0@              &@      $@       @       @              �?       @      �?       @                      �?      @       @              @      @      �?      �?      �?              �?      �?               @              $@       @       @               @       @      �?       @              @      �?      �?      �?                      �?      �?              @      0@      @      @      @               @      @              @       @                      $@      Y@     �u@      A@     `m@      0@      0@       @      ,@       @       @              @       @      �?       @                      �?              @      ,@       @      @      �?      @                      �?      &@      �?      �?      �?      �?                      �?      $@              2@     `k@             �I@      2@      e@       @              0@      e@      (@     `d@      &@     @]@      @     @U@      @     �J@      @      7@      @      @      @      @      @      @      �?      @              @      �?              @                      �?              @              0@              >@              @@      @      @@      @      3@      @      @      @              �?      @              @      �?                      0@              *@      �?      G@              C@      �?       @              @      �?      @              @      �?              @      @              @      @             �P@     �[@     �L@     @R@     �D@      ,@     �C@      &@      <@      &@      @      @              @      @              6@       @      @              0@       @              �?      0@      @      *@      @       @      @       @      @      @      @      @       @       @              �?       @      �?      �?      �?                      �?              �?              �?      @                       @      @       @      @                       @      @              &@               @      @              @       @              0@     �M@      @       @      @                       @      *@     �L@      @     �H@      @     �H@      @      5@      @      $@              "@      @      �?              �?      @                      &@              <@       @              @       @      @       @      @      �?      �?      �?              �?      �?               @              @      �?              �?      @                      @      "@     �B@      @      @              @      @               @      >@       @      (@              &@       @      �?       @                      �?              2@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ/��hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKͅ�h��B@3         T       
             �?4�5����?�           ��@               #                    �?`}�?��?�            �t@,0,Up,0                          �P@���ۑ��?x            �h@      @                           �?և���X�?             ,@     �?                           �?���!pc�?             &@       ������������������������       �                      @      �?������������������������       �                     @        ������������������������       �                     @      �?	                           @L@@-�_ .�?p             g@     �?
                          �g@pY���D�?`            �c@     �?                          @[@ u�z\A�?_            `c@      &@                           @G@�C��2(�?             &@      �?������������������������       �                      @      $@                           �?�q�q�?             @        ������������������������       �                     �?      �?                          `m@      �?              @        ������������������������       �                     �?t,1
54,������������������������       �                     �?        ������������������������       �        Y             b@        ������������������������       �                     @B��fn       "                    �?�<ݚ�?             ;@                                 Pc@���Q��?
             .@                                  �?z�G�z�?             $@                                 �`@�q�q�?             @ �`3���                          @b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     @               !                    �N@z�G�z�?             @                      	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @      C@������������������������       �                      @      @������������������������       �                     (@        $       K                    �?�c��{-�?P            ``@     &@%       0                    �?���I���?A            �[@        &       /                    @d��0u��?             >@     �?'       .                   pf@��X��?             <@     @(       +                   @b@R�}e�.�?             :@      @)       *                   �t@�X�<ݺ?             2@     �?������������������������       �                     1@       @������������������������       �                     �?        ,       -                   �\@      �?              @     �M@������������������������       �                      @     �L@������������������������       �                     @      $@������������������������       �                      @        ������������������������       �                      @       @1       <                   �_@ޭ�W[��?,            @T@      �?2       ;                    _@#z�i��?            �D@     �?3       :       	          ����?4�2%ޑ�?            �A@     @4       9                    ]@ףp=
�?             >@     (@5       6                   �b@z�G�z�?	             .@     �?������������������������       �                     &@        7       8                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     @        ������������������������       �                     @        =       D                   �b@      �?             D@       >       ?                    @M@ >�֕�?            �A@       ������������������������       �                     ;@        @       A                   �c@      �?              @       ������������������������       �                     @        B       C                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        E       J                    @���Q��?             @       F       I       	          `ff�?�q�q�?             @       G       H                    �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        L       S       	          433�?R���Q�?             4@        M       R                   ``@�q�q�?             "@       N       O                    �I@؇���X�?             @       ������������������������       �                     @        P       Q                    ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        U       �                    �?P� �&�?           @y@       V       �                   �b@4��2�?�            u@       W       �                    �R@������?�            �q@       X       �                    @$��{~�?�            �q@       Y       \                   �Q@`q�����?�             q@        Z       [                    Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       �                    �?X�Հ�+�?�            �p@       ^       �                     P@�D����?}            �f@       _       |                   �p@�S(��d�?k            @c@       `       w                   8p@t��%�?U            �\@       a       v                   �m@h�)S;�?Q            �[@       b       k                   `_@�ɮ����?D            �V@       c       h                   �l@h㱪��?+            �K@       d       e                    @O@���J��?'            �I@       ������������������������       �        "            �F@        f       g                    `@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        i       j       	          `ff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        l       q                   �\@tk~X��?             B@        m       p                    �H@      �?             $@       n       o                   �k@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        r       u       	          ����?$�q-�?             :@        s       t                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     3@        x       y                    �K@���Q��?             @        ������������������������       �                     �?        z       {                    @O@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        }       �                    �? ���J��?            �C@        ~                          �`@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@        ������������������������       �                     ;@        �       �                   �`@�x�E~�?2            @V@       ������������������������       �        )            �R@        �       �                    �?�r����?	             .@        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �i@���!pc�?             &@        ������������������������       �                     @        �       �       	          ���@���Q��?             @       �       �                   �j@      �?             @        ������������������������       �                      @        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �[@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    ]@x�K��?            �I@        �       �                    Y@؇���X�?             ,@        ������������������������       �                     @        �       �                   `m@z�G�z�?             $@        ������������������������       �                     @        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        �       �                   `\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��+��?            �B@        �       �       	          `ff@z�G�z�?
             4@       ������������������������       �                     &@        �       �       	          `ff@X�<ݚ�?             "@        ������������������������       �                      @        �       �                   (p@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   pc@�t����?
             1@        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                    �?B�
k���?+            �P@       �       �       	             @�^���U�?$            �L@       �       �                    �?�z�G��?              I@        �       �                   @m@D�n�3�?             3@        ������������������������       �                     @        �       �                    �?d}h���?	             ,@       �       �                   �s@r�q��?             (@       ������������������������       �                     "@        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �g@��� ��?             ?@        �       �                   d@      �?             @       �       �                   @[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �? 7���B�?             ;@       ������������������������       �                     3@        �       �                    �?      �?              @       �       �                   �a@z�G�z�?             @        ������������������������       �                     @        �       �       	          `ff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       �t@     y@     0p@     �Q@     �f@      0@       @      @       @      @       @                      @              @     �e@      $@     @c@      @     @c@      �?      $@      �?       @               @      �?      �?              �?      �?      �?                      �?      b@                      @      5@      @      "@      @       @       @      @       @      �?       @               @      �?              @              @              �?      @      �?       @      �?                       @               @      (@              S@     �K@     @R@      C@      &@      3@      "@      3@      @      3@      �?      1@              1@      �?              @       @               @      @               @               @              O@      3@      ;@      ,@      ;@       @      ;@      @      (@      @      &@              �?      @      �?                      @      .@                      @              @     �A@      @     �@@       @      ;@              @       @      @              �?       @               @      �?               @      @       @      �?      �?      �?              �?      �?              �?                       @      @      1@      @      @      �?      @              @      �?       @      �?                       @       @                      &@     �R@     �t@     �C@     �r@      3@     �p@      2@     �p@      .@     p@      �?      �?              �?      �?              ,@      p@      (@      e@      (@     �a@      &@      Z@      "@     @Y@      "@     �T@       @     �J@      �?      I@             �F@      �?      @      �?                      @      �?      @      �?                      @      @      =@      @      @       @      @              @       @              @               @      8@       @      �?       @                      �?              7@              3@       @      @      �?              �?      @              @      �?              �?      C@      �?      @      �?                      @              @@              ;@       @     �U@             �R@       @      *@       @      @       @                      @               @      @       @              @      @       @      @      �?       @              �?      �?              �?      �?                      �?      �?       @              �?      �?      �?              �?      �?              4@      ?@       @      (@              @       @       @              @       @      �?      �?              �?      �?      �?                      �?      2@      3@      0@      @      &@              @      @               @      @       @      @                       @       @      .@       @      �?       @                      �?              ,@     �A@      @@     �A@      6@     �A@      .@       @      &@      @              @      &@       @      $@              "@       @      �?       @                      �?      �?      �?              �?      �?              ;@      @      �?      @      �?      �?      �?                      �?               @      :@      �?      3@              @      �?      @      �?      @              �?      �?              �?      �?              @                      @              $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJu�7hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKׅ�h��B�5         N       	          ����?p�Vv���?�           ��@      @                           �?X~�pX��?�            �v@               
       
             �?��y�:�?,            �P@      �?                           �B@      �?             @@      �?������������������������       �                     @     �O@                          �h@8^s]e�?             =@      E@������������������������       �                     @      K@       	                     R@�C��2(�?             6@    �N@������������������������       �                     4@Xyrr   r������������������������       �                      @
                            c@ >�֕�?            �A@�              	          ����?г�wY;�?             A@
������������������������       �                     <@      	                            `@r�q��?             @ | dd�������������������������       �                     �? j	t|�������������������������       �                     @the mode������������������������       �                     �?t,1
54,       9       
             �?BA�V�?�            �r@              2                   �b@ d�=��?�            @l@                                  U@X�?٥�?�            �i@ B��fn������������������������       �                     �?              !       	          ����?��?ȿ}�?�            �i@                                  �?����ȫ�?h            �d@       ������������������������       �        P            �_@ �`3���                           d@@-�_ .�?            �B@       ������������������������       �                     <@                                   �E@�<ݚ�?             "@       ������������������������       �                     @                                  ]@�q�q�?             @        ������������������������       �                     �?                                  �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?     �R@"       /                   @n@��r._�?            �D@     @#       (       	          833�?(N:!���?            �A@       @$       %                    �?����X�?             @     �?������������������������       �                     @      �?&       '                    ]@�q�q�?             @      ?@������������������������       �                      @      @������������������������       �                     �?        )       *                    Z@@4և���?             <@        ������������������������       �                     �?        +       ,                    c@ 7���B�?             ;@       ������������������������       �        
             6@      6@-       .                    @F@z�G�z�?             @      &@������������������������       �                     �?        ������������������������       �                     @        0       1                   �_@      �?             @        ������������������������       �                     @        ������������������������       �                     @      �?3       4                   d@�z�G��?             4@      @������������������������       �                     $@        5       8                    �?���Q��?             $@       6       7                   @g@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        :       E                   �b@      �?0             R@       ;       D                   pm@�:�^���?            �F@       <       A                   k@؇���X�?             <@       =       @                    �L@���7�?             6@        >       ?       	          ����?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             *@        B       C                   `^@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             1@        F       M                   0f@|��?���?             ;@       G       H                    �D@�q�q�?             8@        ������������������������       �                     @        I       J                   q@�d�����?             3@       ������������������������       �                     *@        K       L                    @O@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        O       �                   �b@�zц��?�            w@       P       _       
             �?+FJ�?�            �r@        Q       Z                    @L@H�z�G�?             D@        R       Y                    �?�d�����?
             3@        S       X       	             �?      �?              @       T       W                    �?���Q��?             @        U       V                   @a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        [       \                    c@؇���X�?             5@       ������������������������       �                     1@        ]       ^                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        `       s                    �?������?�            0p@        a       r                   �s@      �?             D@       b       k                   pa@�θ�?            �C@       c       d                   l@�����H�?             2@       ������������������������       �        	             (@        e       f                   �l@�q�q�?             @        ������������������������       �                     �?        g       j                    @K@z�G�z�?             @        h       i                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        l       q                   o@�q�q�?             5@        m       p       	          `ff@�<ݚ�?             "@       n       o                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        t       �                   `\@ �o�b��?�            `k@        u       �                    @Q@�<ݚ�?             B@       v       �                    �?      �?             @@       w       x                   `_@8�Z$���?             :@        ������������������������       �        	             &@        y       �                   �b@������?
             .@       z       �                   0b@�q�q�?             (@       {       �                    �?z�G�z�?             $@       |       �                   �a@�<ݚ�?             "@       }       �                   �m@�q�q�?             @       ~                            E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �L@�]0��<�?z            �f@       �       �                    �?�X�<ݺ??            �V@       �       �       	          ����?(�5�f��?6            �S@        �       �       	          `ff�?r�q��?             (@        ������������������������       �                     @        �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        �       �                   @[@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          033@�\=lf�?.            �P@       ������������������������       �        $             K@        �       �                   �\@$�q-�?
             *@        �       �                    �J@      �?             @        �       �                    @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   @[@"pc�
�?	             &@        ������������������������       �                     @        �       �                   �p@      �?              @        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `\@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�L��ȕ?;            @W@       ������������������������       �        ,            @R@        �       �                    `@P���Q�?             4@        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        �       �                    �?��(@��?.            �Q@       �       �                    �L@�eP*L��?"            �K@       �       �                    �?�q�q�?            �@@       �       �                    U@\X��t�?             7@        ������������������������       �                     @        �       �       
             �?��Q��?             4@       �       �       	             @�E��ӭ�?             2@       �       �                   pc@     ��?
             0@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �G@$�q-�?             *@       ������������������������       �                      @        �       �                   0`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?ףp=
�?             $@        �       �       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pc@���|���?             6@        �       �                    �O@      �?              @        �       �       	          033�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �c@@4և���?	             ,@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �d@z�G�z�?             .@        �       �                     K@      �?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @       �       �                   �c@      �?             @        ������������������������       �                     �?        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �t�bh�h*h-K ��h/��R�(KK�KK��ha�Bp       @t@     �y@     @o@     �\@      6@     �F@      4@      (@              @      4@      "@              @      4@       @      4@                       @       @     �@@      �?     �@@              <@      �?      @      �?                      @      �?             �l@     �Q@     @j@      0@     �h@      $@              �?     �h@      "@     @d@       @     �_@             �A@       @      <@              @       @      @              �?       @              �?      �?      �?              �?      �?              A@      @      ?@      @      @       @      @              �?       @               @      �?              :@       @              �?      :@      �?      6@              @      �?              �?      @              @      @              @      @              ,@      @      $@              @      @      @      �?      @                      �?              @      2@      K@      @     �D@      @      8@      �?      5@      �?       @               @      �?                      *@      @      @              @      @                      1@      ,@      *@      ,@      $@              @      ,@      @      *@              �?      @              @      �?                      @     �R@     pr@     �D@      p@      1@      7@      ,@      @      @      @      @       @      �?       @               @      �?               @                      @      &@              @      2@              1@      @      �?      @                      �?      8@     `m@      $@      >@      "@      >@       @      0@              (@       @      @      �?              �?      @      �?      �?              �?      �?                      @      @      ,@      @       @      @      �?              �?      @                      �?              (@      �?              ,@     �i@       @      <@      @      <@      @      6@              &@      @      &@      @       @       @       @       @      @       @      @       @      �?              �?       @                      @              @              �?       @                      @              @      @              @      f@      @     @U@      @      S@       @      $@              @       @      @               @       @      @       @                      @      �?     �P@              K@      �?      (@      �?      @      �?      �?              �?      �?                       @              "@       @      "@              @       @      @      �?      �?      �?                      �?      �?      @      �?                      @      �?      W@             @R@      �?      3@      �?      �?              �?      �?                      2@     �@@     �B@      >@      9@      6@      &@      *@      $@              @      *@      @      *@      @      *@      @      �?       @      �?                       @      (@      �?       @              @      �?              �?      @                       @               @      "@      �?       @      �?       @                      �?      @               @      ,@      @      �?      @      �?              �?      @              @              �?      *@      �?      @              @      �?                      $@      @      (@      @      @              �?      @       @       @       @              �?       @      �?              �?       @              �?                      "@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��!XhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B@/         N                    �?U�ք�?�           ��@      (@       K                    @JN�#:�?�            �s@,180,0,              
             �?��A�J��?�            0s@     �@@                           I@�p ��?            �D@      @                           `@�C��2(�?             &@      @������������������������       �                     $@       @������������������������       �                     �?      �?              	          ����?�q�q�?             >@       	                            R@��s����?             5@       
                           �I@�KM�]�?             3@       ������������������������       �                     $@                                   �?�<ݚ�?             "@       ������������������������       �                     @                                  �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                  �`@�q�q�?             "@     @                          �^@      �?             @      @������������������������       �                      @      p@                          �r@      �?             @      @������������������������       �                     @        ������������������������       �                     �?      1@������������������������       �                     @     `m@       :                    a@��i��X�?�            �p@     (@              	          ����?8be��|�?             i@      �?������������������������       �                     =@      ,@       /                    \@�Ts�k��?k            �e@               .                    @R@�t����?)             Q@    �i@              	          hff�?$�q-�?(            @P@      &@������������������������       �                     �?      @        !                    h@      �?'             P@        ������������������������       �                     6@        "       -                    �L@�����?             E@     f@#       $                   Pj@�㙢�c�?             7@      @������������������������       �                     �?        %       &                    �H@��2(&�?             6@      (@������������������������       �                     $@        '       (                    �I@      �?             (@      @������������������������       �                     �?      �?)       *                   �Z@"pc�
�?             &@     W@������������������������       �                      @      �?+       ,       	          033@�q�q�?             @     9@������������������������       �                      @      @������������������������       �                     �?        ������������������������       �                     3@      �?������������������������       �                     @       @0       9                   P`@��9J���?B             Z@      �?1       8                   �_@t��ճC�?             F@     �?2       3                    @L@ �Cc}�?             <@     *@������������������������       �                     2@      $@4       7                    �N@�z�G��?             $@      @5       6                   �d@      �?             @      �?������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �        #             N@        ;       J                   pn@؇>���?*            @P@       <       G                    �?��J�fj�?            �B@       =       F                    �?���Q��?             9@       >       A                    `@�\��N��?             3@        ?       @                   `h@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        B       C                   `d@z�G�z�?             $@       ������������������������       �                     @        D       E                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        H       I                   Pa@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     <@        L       M                    �C@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        O       |       
             �?n�����?           @z@       P       [                   @E@����y7�?�            @o@        Q       X                   P`@�q�q�?             2@       R       W                    �?8�Z$���?
             *@        S       T                    �?�q�q�?             @        ������������������������       �                     �?        U       V       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        Y       Z                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        \       u                    �O@�8���?�             m@       ]       t                   h@�v�ɱ?�            �k@       ^       s       	          ���@p���4h�?�            �k@       _       j                   Pb@Ц�f*�?�            �k@       `       a                    �?     ��?}             h@       ������������������������       �        h            @d@        b       e                    @F@ףp=
�?             >@        c       d                    �?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        f       g                    �?�}�+r��?             3@       ������������������������       �                     0@        h       i                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        k       l                    �? �Cc}�?             <@       ������������������������       �                     5@        m       r                   Hq@և���X�?             @       n       o                   �d@      �?             @        ������������������������       �                      @        p       q                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        v       {                    �P@���Q��?             $@       w       x                    ]@      �?              @        ������������������������       �                      @        y       z       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        }       �                    �?f��>���?o            @e@       ~       �                   c@6YE�t�?U            �`@              �                    �?�^'�ë�?=            @X@       �       �       	          ����?��}���?3            @S@        ������������������������       �                     <@        �       �                   �]@�����?            �H@        �       �                    �M@�IєX�?
             1@        �       �       	             �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?     ��?             @@       �       �       	          033�?�G�z��?             4@        ������������������������       �                     @        �       �       
             �?d}h���?             ,@       �       �       	          ����?�8��8��?             (@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �        
             4@        �       �       	             @����X�?            �A@       �       �                   �i@r٣����?            �@@        ������������������������       �                     $@        �       �                   `\@�LQ�1	�?             7@        ������������������������       �                     @        �       �                   0f@���Q��?             4@       �       �                   `]@�q�q�?             2@        ������������������������       �                      @        �       �       	          `ff�?      �?             0@       �       �       
             �?����X�?
             ,@       �       �                   0`@�θ�?	             *@        ������������������������       �                     @        �       �       	          hff�?�q�q�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        �       �                   0m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �       	          ��� @D�n�3�?             C@       �       �                    `P@�4�����?             ?@       �       �                    @N@���Q��?             9@       �       �                   �Q@      �?             4@        ������������������������       �                      @        �       �                   �b@r�q��?             2@       �       �                    �?�t����?             1@       ������������������������       �                     &@        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     P@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B�        t@     �y@      K@     @p@      H@     0p@      5@      4@      �?      $@              $@      �?              4@      $@      1@      @      1@       @      $@              @       @      @              �?       @      �?                       @               @      @      @      @      @               @      @      �?      @                      �?              @      ;@     �m@      &@     �g@              =@      &@      d@       @      N@      @      N@      �?              @      N@              6@      @      C@      @      3@      �?              @      3@              $@      @      "@      �?               @      "@               @       @      �?       @                      �?              3@      @              @     @Y@      @     �D@      @      9@              2@      @      @      @      @              @      @                      @              0@              N@      0@     �H@      0@      5@      .@      $@      "@      $@      @       @               @      @               @       @              @       @      �?              �?       @              @              �?      &@      �?                      &@              <@      @      �?              �?      @             �p@      c@     @l@      8@      @      (@       @      &@       @      �?      �?              �?      �?      �?                      �?              $@      @      �?      @                      �?     �k@      (@     �j@       @     �j@      @     �j@      @     �g@      @     @d@              ;@      @      "@       @      "@                       @      2@      �?      0@               @      �?       @                      �?      9@      @      5@              @      @      �?      @               @      �?      �?              �?      �?              @                      �?              �?      @      @      @      @               @      @       @               @      @               @              E@      `@      4@      \@      $@     �U@      $@     �P@              <@      $@     �C@      �?      0@      �?      @      �?                      @              $@      "@      7@      "@      &@      @              @      &@      �?      &@      �?       @      �?                       @              "@       @                      (@              4@      $@      9@       @      9@              $@       @      .@              @       @      (@      @      (@               @      @      $@      @      $@      @      $@              @      @      @              @      @      @      �?       @               @      �?               @      �?       @                      �?      �?               @               @               @              6@      0@      5@      $@      .@      $@      .@      @               @      .@      @      .@       @      &@              @       @      @                       @              �?              @      @              �?      @              @      �?        �t�bub�     hhubh)��}�(hhhhhNhKhKhG        hh&hNhJC�NhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK�h��B@<         V                    �?4�5����?�           ��@      �?                           �?Z�/�j��?�            �r@ ,ATA,12                           �?��N`.�?'            �K@       @              
             �?
j*D>�?             :@       @������������������������       �                     "@                                  `f@ҳ�wY;�?             1@        ������������������������       �                     @               	                    �J@      �?	             (@        ������������������������       �                     @        
                          s@؇���X�?             @       ������������������������       �                     @                                  xt@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?ܷ��?��?             =@       ������������������������       �                     9@                                  @_@      �?             @ �s��  ������������������������       �                      @given RV                           �?      �?              @ y_like
������������������������       �                     �?ay_like
������������������������       �                     �?(see doc       !                   �]@T$�#���?�            `n@ ation)
                           `@X�<ݚ�?             2@ aramete                           �?      �?              @      s              	          �����      �?             @ --
    ������������������������       �                     �?on evalu������������������������       �                     @ r   r�������������������������       �                     @ r   �                           �?ףp=
�?             $@r�   r�������������������������       �                     @  s"                             @b@      �?             @        ������������������������       �                     @}}tt������������������������       �                     �?      @"       M       	          033�?��1�'��?�             l@     7@#       2       
             �?0��_��?�            �j@     &@$       /                    �?`<�Gf�?r             e@     "@%       .                   �c@@��t��?a             b@     9@&       -                   xt@hA� �?2            �Q@     @'       ,                    �G@ ��ʻ��?1             Q@      $@(       +                    �?�g�y��?             ?@     @)       *                   �\@ �q�q�?             8@       @������������������������       �                     �?      �?������������������������       �                     7@        ������������������������       �                     @      @������������������������       �                    �B@        ������������������������       �                      @      �?������������������������       �        /            �R@      @0       1                    f@�8��8��?             8@       ������������������������       �                     6@        ������������������������       �                      @        3       J                   0a@8�$�>�?            �E@       4       ;                   �a@������?             A@        5       8                    �?�q�q�?             @        6       7                    a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        9       :                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        <       A                   �d@؇���X�?             <@       =       @                    �?���N8�?
             5@        >       ?                    �K@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        B       C                   e@և���X�?             @        ������������������������       �                      @8 +�&� D       I                    �?z�G�z�?             @       E       F                   `\@�q�q�?             @        ������������������������       �                     �?        G       H                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        K       L                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        N       U       	             @�	j*D�?	             *@       O       T                   �r@      �?              @       P       S                    �L@�q�q�?             @       Q       R                   pc@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        W       �       	          ����?      �?           @{@        X       k                    �?\`*�s�?k             e@        Y       h                    �?t�F�}�?            �I@       Z       [                    �F@^H���+�?            �B@        ������������������������       �                     @        \       ]                   �_@*;L]n�?             >@        ������������������������       �                     $@        ^       e                    �?��Q��?             4@       _       `       
             �?և���X�?
             ,@        ������������������������       �                     @        a       d                   �\@�q�q�?             "@        b       c                    Y@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        f       g                   �\@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        i       j                    @J@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        l       �                    �?z4��f��?L            @]@       m       |                   `_@ƈ�VM�?:            @V@        n       u                    �?*;L]n�?             >@        o       t                   `c@؇���X�?             ,@       p       s                    @I@$�q-�?             *@        q       r                   @Z@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        v       {       	          @33�?     ��?             0@       w       x                   @\@�8��8��?             (@       ������������������������       �                     @        y       z       
             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        }       �       
             �?L
�q��?*            �M@       ~       �       	            �?���?            �D@              �                    @F@x�����?            �C@        �       �                   `i@ҳ�wY;�?             1@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �e@r�q��?	             (@       �       �                    �?�C��2(�?             &@       �       �                    �E@ףp=
�?             $@       ������������������������       �                      @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    s@�C��2(�?             6@       �       �                    @N@���N8�?             5@       ������������������������       �                     .@        �       �                    �N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �_@X�<ݚ�?             2@        ������������������������       �                     @        �       �                   0a@���!pc�?             &@        ������������������������       �                     @        �       �                    �N@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?      �?             <@       ������������������������       �                     2@        �       �                   `\@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?��v����?�            �p@        �       �       	          033�?h+�v:�?             A@       �       �                    �?l��
I��?             ;@       �       �                    �?��<b���?             7@       �       �                     F@ףp=
�?             4@        ������������������������       �                     �?        �       �                    c@�}�+r��?             3@       ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �h@����X�?             @        ������������������������       �                     @        �       �       	          033@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @f@�q�6m��?�            @m@       �       �                   �Q@��Q�Vz�?�            �l@        �       �                    �N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?0�֋���?�            @l@       �       �                   i@@-�_ .�?|             g@        ������������������������       �        *             N@        �       �       	          ����?HP�s��?R            @_@        �       �                   �[@�q�q�?             8@        �       �                   �`@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�S����?             3@       ������������������������       �        
             *@        �       �                   @\@      �?             @       �       �                   @^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   pb@��^M}�?B            @Y@       �       �                    _@�g�y��?:            @W@        �       �                   Pk@�r����?             .@        ������������������������       �                     �?        �       �       	          ���@@4և���?
             ,@       ������������������������       �                     "@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   Ps@�(�Tw�?/            �S@       ������������������������       �        $            �M@        �       �                    �?�}�+r��?             3@       ������������������������       �        
             2@        ������������������������       �                     �?        �       �                    \@      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @       �       �                    q@      �?             @        ������������������������       �                      @        �       �                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��r._�?            �D@       �       �                   h@�'�`d�?            �@@        �       �                   �R@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `P@\-��p�?             =@       �       �                   �q@ �Cc}�?             <@        ������������������������       �                     1@        �       �       	          ����?���!pc�?             &@        �       �                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `]@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B       �t@     y@      l@     �R@      2@     �B@      .@      &@      "@              @      &@              @      @      @      @              �?      @              @      �?       @      �?                       @      @      :@              9@      @      �?       @              �?      �?              �?      �?             �i@     �B@      $@       @      �?      @      �?      @      �?                      @              @      "@      �?      @              @      �?      @                      �?     �h@      =@      h@      4@     �d@      @     �a@      @     �P@      @     �P@      �?      >@      �?      7@      �?              �?      7@              @             �B@                       @     �R@              6@       @      6@                       @      <@      .@      :@       @       @      @      �?      @      �?                      @      �?      �?              �?      �?              8@      @      4@      �?      @      �?      @                      �?      ,@              @      @               @      @      �?       @      �?      �?              �?      �?      �?                      �?       @               @      @              @       @              @      "@      @      @       @      @       @      �?              �?       @                      @       @                      @     @[@     pt@     @R@     �W@      ,@     �B@      *@      8@              @      *@      1@              $@      *@      @       @      @      @              @      @      @      �?              �?      @                      @      @      �?              �?      @              �?      *@      �?                      *@     �M@      M@      J@     �B@      *@      1@       @      (@      �?      (@      �?      @      �?                      @              @      �?              &@      @      &@      �?      @              @      �?      @                      �?              @     �C@      4@      ?@      $@      ?@       @      &@      @      �?      @              @      �?              $@       @      $@      �?      "@      �?       @              �?      �?      �?                      �?      �?                      �?      4@       @      4@      �?      .@              @      �?              �?      @                      �?               @       @      $@              @       @      @      @               @      @              @       @              @      5@              2@      @      @              @      @              B@      m@      *@      5@       @      3@      @      2@       @      2@      �?              �?      2@              2@      �?              @              @      �?      �?      �?              �?      �?               @              @       @      @              �?       @      �?                       @      7@     `j@      3@     @j@       @      �?       @                      �?      1@      j@      $@     �e@              N@      $@     �\@      @      3@       @      @              @       @              @      0@              *@      @      @      @      �?              �?      @                       @      @      X@      @     �V@       @      *@      �?              �?      *@              "@      �?      @              @      �?              �?     @S@             �M@      �?      2@              2@      �?               @      @      �?              �?      @      �?      @               @      �?      �?      �?                      �?              @      @      A@      @      :@      @      �?              �?      @              @      9@      @      9@              1@      @       @      @      �?      @                      �?              @      �?                       @      @      �?      @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�R�[hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKۅ�h��B�6         `       	          ����?6������?�           ��@              E       
             �?��_���?�             w@,N,1,Fl                          @E@(��R%��?�            �p@       @                          �[@��H�}�?             9@      9@������������������������       �                     @     �G@                           �?�\��N��?             3@     F@                           �?���Q��?	             .@    �I@                           �?      �?             (@     �G@	       
                   �a@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?                                  @_@�����H�?             "@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                     @        ������������������������       �                     @      �?������������������������       �                     @               6                   q@�l�T{�?�             n@     @       3       	          ����?�g��.��?v            �f@     @                          �b@�ȨF=�?t            `f@     @                          �a@�����??            @Y@    �W@������������������������       �        *             Q@      1@                          p@Pa�	�?            �@@       ������������������������       �                     ?@                                   �H@      �?              @        ������������������������       �                     �?      M@������������������������       �                     �?      (@       ,                    @M@$�q-�?5            �S@     @       )                   �b@�X�<ݺ?1             R@              "                   �e@��.N"Ҭ?/            @Q@      @        !                   �\@ףp=
�?             $@      @������������������������       �                     �?       @������������������������       �                     "@      �?#       (                   @[@P����?)            �M@      �?$       '                    �?r�q��?             @      �?%       &                    c@      �?              @       @������������������������       �                     �?        ������������������������       �                     �?      5@������������������������       �                     @        ������������������������       �        %            �J@      2@*       +                   �c@�q�q�?             @      2@������������������������       �                      @      �?������������������������       �                     �?       @-       .                   �`@�q�q�?             @       @������������������������       �                     @        /       2                    b@�q�q�?             @     N@0       1                    �?      �?              @      @������������������������       �                     �?      @������������������������       �                     �?       @������������������������       �                     �?        4       5                   p@      �?              @      @������������������������       �                     �?      2@������������������������       �                     �?        7       >                    �L@z�G�z�?&             N@     �?8       9                    �?�����?             E@     A@������������������������       �                    �A@        :       =                    @F@և���X�?             @      @;       <                   �r@z�G�z�?             @     @������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ?       D                    �?X�<ݚ�?             2@       @       A                   �c@�C��2(�?             &@       ������������������������       �                      @        B       C                   @`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        F       S       	          ����?�4�M�f�?@            �Y@       G       H                   Pi@86��Z�?0            �S@       ������������������������       �                     D@        I       R                   0a@�ݜ�?            �C@       J       O                    �?z�G�z�?             9@       K       N       
             �?؇���X�?             5@       L       M                   �i@�}�+r��?
             3@        ������������������������       �                     �?        ������������������������       �        	             2@        ������������������������       �                      @        P       Q                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        T       U                   �g@�û��|�?             7@        ������������������������       �                     @        V       Y                    �?�d�����?             3@        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       _                   �q@     ��?	             0@       [       ^                    `@@4և���?             ,@        \       ]                   `o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        a       �                   �`@xƅd�?�            �v@       b       g                    �?ܷ��?��?~            `i@        c       f                   Pm@      �?             @       d       e       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        h       �                    �Q@�����?z            �h@       i       �       
             �?��Y���?u            �g@       j       y                   �_@0��P�?g            �d@        k       l                   `[@��0{9�?            �G@        ������������������������       �                     0@        m       n                   �h@��a�n`�?             ?@        ������������������������       �                     *@        o       p                   �\@b�2�tk�?             2@        ������������������������       �                     @        q       v                    �K@d}h���?
             ,@       r       s                    _@�����H�?             "@       ������������������������       �                     @        t       u       	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        w       x                    @M@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        z       �                    `@ ���J��?L            @]@       {       �                   P`@���1��?C            �Z@        |       }                    �?      �?             0@       ������������������������       �                     *@        ~                           �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        ;            �V@        �       �       
             �?z�G�z�?	             $@        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @       ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                   Xs@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   (w@�+$�jP�?             ;@       �       �                    �?H%u��?             9@       ������������������������       �        	             0@        �       �                   �]@�q�q�?             "@       �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?噼:��?d            `d@        �       �       	          ����?      �?-             R@        �       �                   �m@ףp=
�?             4@       ������������������������       �                     ,@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �k@�	j*D�?              J@        �       �                    �?�q�q�?             8@        ������������������������       �                      @        �       �       	          033�?      �?             0@        ������������������������       �                     �?        �       �                    �?�q�q�?             .@       �       �                    @I@r�q��?	             (@        ������������������������       �                     @        �       �       
             �?      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @       �       �                   �X@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    a@@4և���?             <@        ������������������������       �                     .@        �       �                    �?8�Z$���?	             *@        �       �                   �b@����X�?             @        ������������������������       �                     @        �       �                   pd@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @L@fK!���?7            �V@       �       �       	          033@ �o_��?             I@       �       �                    �?r�q��?             E@       �       �                   `U@R�}e�.�?             :@        ������������������������       �                      @        �       �       
             �?�q�q�?             8@       �       �                    a@��2(&�?             6@       �       �                   �a@�X�<ݺ?             2@        �       �       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             .@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             0@        �       �       
             �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   `a@���� �?            �D@        ������������������������       �                      @        �       �       	          ����?�θ�?            �C@        �       �                    �?�eP*L��?             &@       �       �                   n@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? �Cc}�?             <@        �       �                   �_@�q�q�?             "@       ������������������������       �                     @        �       �       	          ���@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             3@        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       �t@     �x@      o@     �]@     �l@      B@      "@      0@              @      "@      $@      "@      @      "@      @      �?       @               @      �?               @      �?       @      �?              �?       @              @                      @              @     �k@      4@     �e@       @     �e@      @      Y@      �?      Q@              @@      �?      ?@              �?      �?      �?                      �?      R@      @      Q@      @     �P@       @      "@      �?              �?      "@              M@      �?      @      �?      �?      �?              �?      �?              @             �J@              �?       @               @      �?              @       @      @              �?       @      �?      �?      �?                      �?              �?      �?      �?              �?      �?              H@      (@      C@      @     �A@              @      @      �?      @              @      �?               @              $@       @      $@      �?       @               @      �?       @                      �?              @      3@     �T@      @     �R@              D@      @      A@      @      4@      @      2@      �?      2@      �?                      2@       @               @       @       @                       @              ,@      ,@      "@              @      ,@      @      �?       @      �?                       @      *@      @      *@      �?      �?      �?              �?      �?              (@                       @     �U@     �q@      5@     �f@       @       @       @      �?              �?       @                      �?      3@     �f@      .@      f@      $@     @c@      @      D@              0@      @      8@              *@      @      &@      @              @      &@      �?       @              @      �?       @      �?                       @       @      @       @                      @      @     �\@      �?     �Z@      �?      .@              *@      �?       @      �?                       @             �V@       @       @      �?      �?      �?                      �?      �?      @              @      �?       @      �?      �?      �?                      �?              �?      @      6@      @      6@              0@      @      @      �?      @      �?                      @       @               @              @      @      @                      @     @P@     �X@      2@      K@       @      2@              ,@       @      @       @                      @      0@      B@      ,@      $@       @              @      $@      �?              @      $@       @      $@              @       @      @      �?              �?      @      �?      @      �?                      @              @      @               @      :@              .@       @      &@       @      @              @       @      �?       @                      �?              @     �G@      F@      B@      ,@     �A@      @      3@      @               @      3@      @      3@      @      1@      �?       @      �?       @                      �?      .@               @       @       @                       @               @      0@              �?      @              @      �?              &@      >@       @              "@      >@      @      @      �?      @              @      �?              @              @      9@      @      @              @      @      �?      @                      �?              3@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�v}hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK݅�h��B@7         f                    �?U�ք�?�           ��@      0@       9                    @L@������?�            �r@              
                    I@ޗQ�~�?�            �i@      �?                           @J@�q�q�?             (@                     	          �����؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @      �?       	                    �?z�G�z�?             @        ������������������������       �                     @     �?������������������������       �                     �?     �?       6                   h@      �?             h@     &@       #       	          ����?p�/E�f�?}            �g@     �?                           �?�%IM��?c            �a@     $@                           �?�E�����?=            �V@                                  �? �)���?8            @T@     �?                           �B@�h����?&             L@                      
             �?ףp=
�?	             $@     �?������������������������       �                     "@      D@������������������������       �                     �?      2@������������������������       �                     G@       @������������������������       �                     9@      "@������������������������       �                     "@                      
             �?@�0�!��?&            �I@     �?                           �G@Du9iH��?             �E@       @                          0n@؇���X�?             5@     �?������������������������       �                     ,@     �f@                          @c@և���X�?             @      0@������������������������       �                     @        ������������������������       �                     @       @������������������������       �                     6@               "       	             �?      �?              @     .@        !                   �l@؇���X�?             @       @������������������������       �                     �?        ������������������������       �                     @       @������������������������       �                     �?      �?$       %       
             �?��|�5��?            �G@      @������������������������       �                     ,@        &       '                   @[@�q�q�?            �@@      @������������������������       �                      @      ,@(       3                    �?f���M�?             ?@     B@)       .                    �G@�eP*L��?             6@        *       +       	             @ףp=
�?             $@     @������������������������       �                      @        ,       -                    �?      �?              @      :@������������������������       �                     �?      @������������������������       �                     �?      @/       0       	          ����?      �?             (@     @������������������������       �                     @      �?1       2                    �?���Q��?             @        ������������������������       �                      @       @������������������������       �                     @        4       5                    �K@�����H�?             "@     @������������������������       �                      @        ������������������������       �                     �?      �?7       8                    d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        :       K                    �?�q�q��?:             X@        ;       @                   �m@���y4F�?             C@        <       =       	          033�?P���Q�?             4@       ������������������������       �        	             2@        >       ?                    c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        A       B       
             �?b�2�tk�?             2@        ������������������������       �                     @        C       D                   �n@d}h���?	             ,@        ������������������������       �                      @        E       F                   �s@�8��8��?             (@       ������������������������       �                      @        G       J                    �?      �?             @       H       I                   @[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        L       S                    U@T����1�?$             M@        M       N                   @]@      �?              @        ������������������������       �                     �?        O       P                   �b@؇���X�?             @       ������������������������       �                     @        Q       R                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       a                    �?�-���?             I@       U       \       
             �?����"�?             =@        V       [                    �?��S�ۿ?	             .@        W       X                   Hp@      �?              @        ������������������������       �                     @        Y       Z                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ]       ^                   �a@����X�?
             ,@        ������������������������       �                     @        _       `                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        b       e                   �Z@�����?             5@        c       d       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             2@        g       �       	          ����?Ƶ�pD�?            {@        h       o                    P@�ģ�a@�?j            @e@        i       n                   �Z@г�wY;�?             A@        j       k       	          ���ܿ      �?             @        ������������������������       �                     �?        l       m                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     >@        p       �       	          ����?�hJ,��?Q             a@       q       �                    �?<�;�OK�??            @Y@       r       �                    �L@�G�z�?0             T@       s       �                    @I@���e��?'            �P@       t       �                   �f@�q����?            �J@       u       v                   �a@ \� ���?            �H@        ������������������������       �                      @        w       z                   �a@��[�p�?            �G@        x       y       
             �?b�2�tk�?             2@        ������������������������       �                     @        ������������������������       �                     &@        {       �                    �E@ܷ��?��?             =@       |       �       
             �?@�0�!��?             1@       }       �                    �D@և���X�?             @       ~                          `d@z�G�z�?             @        ������������������������       �                     @        �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     (@        ������������������������       �                     @        �       �       
             �?�	j*D�?	             *@       ������������������������       �                     "@        ������������������������       �                     @        �       �                   �e@@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �J@��s����?             5@       ������������������������       �                     &@        �       �       
             �?���Q��?             $@       �       �                    �N@      �?              @        �       �                    d@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?z�G�z�?            �A@        �       �                    �?�q�q�?             "@       �       �       
             �?���Q��?             @        ������������������������       �                      @        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	            �? ��WV�?             :@       �       �       
             �?      �?             0@       ������������������������       �                     *@        �       �                    b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   P`@�Ra����?�            �p@       �       �                    �R@�;Y�&��?h            @f@       �       �                    �?�f"Nf�?g             f@       �       �                   �]@�(�Tw�?[            �c@       ������������������������       �        :            @Y@        �       �       
             �?h㱪��?!            �K@       �       �                    �?p���?             I@       �       �                   �\@Pa�	�?            �@@        �       �                    @M@      �?             @        �       �                   �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                     1@        �       �       	              @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @����X�?             5@       �       �       	             �?r�q��?
             2@        �       �                   0n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                     �?        �       �                   0i@�������?;            �U@        �       �                   @e@      �?             >@       �       �                    �?8�A�0��?             6@       �       �                     G@���Q��?             .@        ������������������������       �                     @        �       �                    @"pc�
�?             &@       �       �       	             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @      �?              @        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    ]@ �Cc}�?'             L@        �       �                   �a@���Q��?	             $@       �       �                    �I@؇���X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   `a@�nkK�?             G@        ������������������������       �                     3@        �       �                    �?�>����?             ;@       ������������������������       �                     7@        �       �       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B�        t@     �y@     �k@      T@     �e@      ?@      @      @      �?      @      �?                      @      @      �?      @                      �?      e@      8@     �d@      5@     ``@      $@     @V@      �?      T@      �?     �K@      �?      "@      �?      "@                      �?      G@              9@              "@              E@      "@      D@      @      2@      @      ,@              @      @              @      @              6@               @      @      �?      @      �?                      @      �?              B@      &@      ,@              6@      &@       @              4@      &@      (@      $@      "@      �?       @              �?      �?              �?      �?              @      "@              @      @       @               @      @               @      �?       @                      �?      �?      @      �?                      @     �G@     �H@       @      >@      �?      3@              2@      �?      �?              �?      �?              @      &@      @              @      &@       @              �?      &@               @      �?      @      �?      �?              �?      �?                       @     �C@      3@       @      @      �?              �?      @              @      �?      �?              �?      �?             �B@      *@      2@      &@      ,@      �?      @      �?      @              �?      �?              �?      �?              @              @      $@              @      @      @      @                      @      3@       @      �?       @      �?                       @      2@             �Y@     �t@      R@     �X@      �?     �@@      �?      @              �?      �?       @      �?                       @              >@     �Q@     @P@     �E@      M@      :@      K@      9@     �D@      0@     �B@      (@     �B@       @              $@     �B@      @      &@      @                      &@      @      :@      @      ,@      @      @      �?      @              @      �?      �?      �?                      �?       @                      $@              (@      @              "@      @      "@                      @      �?      *@      �?                      *@      1@      @      &@              @      @      @       @       @       @       @                       @      @                       @      <@      @      @      @      @       @       @              �?       @      �?                       @              @      9@      �?      .@      �?      *@               @      �?       @                      �?      $@              >@     @m@      "@      e@       @      e@       @     @c@             @Y@       @     �J@      �?     �H@      �?      @@      �?      @      �?      �?      �?                      �?               @              =@              1@      �?      @      �?                      @      @      .@      @      .@      @      �?              �?      @                      ,@      @              �?              5@     @P@      .@      .@      "@      *@      "@      @              @      "@       @      "@      �?              �?      "@                      �?              @      @       @      �?       @      �?                       @      @              @      I@      @      @      �?      @      �?       @               @      �?                      @      @               @      F@              3@       @      9@              7@       @       @       @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJg}�XhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK�h��B�<         Z                    �?0����?�           ��@                      
             �?�q�� �?�            �r@ 31,0,ST              	          hff�?�Q����?             D@     5@                          0a@     ��?             0@      �?                          �^@����X�?             @        ������������������������       �                     �?      �?       
                   �l@r�q��?             @               	                   �Y@�q�q�?             @        ������������������������       �                      @     �?������������������������       �                     �?     �?������������������������       �                     @     &@������������������������       �                     "@     �?                           c@�q�q�?             8@     $@                          �`@z�G�z�?             4@                                  �^@z�G�z�?             @      �?������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@      �?������������������������       �                     @      3@       9       	          ����?�����?�             p@      @       4                   �b@��k=.��?<            �W@     *@                           �?��|���?8             V@                                   �?�E��ӭ�?             2@                                   @K@X�<ݚ�?             "@        ������������������������       �                     @                                  @_@r�q��?             @     �X@������������������������       �                     �?       @������������������������       �                     @     @P@������������������������       �                     "@     �B@              	          hff�?(N:!���?,            �Q@      &@������������������������       �                     2@      ,@        3                   �a@8�Z$���?!             J@     �?!       "                    �F@���y4F�?             C@      $@������������������������       �                     $@        #       *                   @Z@����X�?             <@      *@$       %                    �?�����H�?             "@       @������������������������       �                     @        &       '                   �Y@z�G�z�?             @       @������������������������       �                      @       @(       )                   (q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @     @c@+       ,                   �i@p�ݯ��?             3@      @@������������������������       �                      @      �?-       .                   �^@���|���?             &@      @������������������������       �                     @      .@/       0                   �`@�q�q�?             @      ,@������������������������       �                     @      .@1       2                   @_@�q�q�?             @       @������������������������       �                      @      �?������������������������       �                     �?        ������������������������       �        	             ,@      @5       6                    �?r�q��?             @        ������������������������       �                     @      3@7       8                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        :       M                   �l@0��P�?g            �d@        ;       F       	          ����?�����?1            �R@        <       E                   0l@z�G�z�?             4@       =       D                    �?�����H�?             2@       >       ?                   �d@�IєX�?             1@       ������������������������       �                     &@        @       C                    �L@r�q��?             @        A       B                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        G       H                   �Z@�X�<ݺ?"             K@        ������������������������       �                      @        I       L                    �? pƵHP�?!             J@        J       K                    [@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     H@        N       W       
             �?(;L]n�?6            �V@       O       V                    c@��Y��]�?0            �T@       P       U                   �_@ �)���?/            @T@        Q       T                   �\@      �?             0@        R       S                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �        $            @P@        ������������������������       �                     �?        X       Y                    �R@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        [       v                   `\@�ua��?           @{@        \       e                   �S@ 1_#�?%            �M@        ]       ^                     G@�8��8��?             8@        ������������������������       �                     �?        _       d       	          ����?�nkK�?             7@       `       a                   �_@      �?             0@       ������������������������       �                     (@        b       c       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        f       u                     P@�xGZ���?            �A@       g       t       	          ����?��S���?             >@       h       m                    �?���!pc�?             6@       i       j                   @Z@؇���X�?
             ,@        ������������������������       �                     @        k       l                   �i@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        n       s                    �?      �?              @       o       p       	             �?�q�q�?             @        ������������������������       �                     @        q       r                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        w       �       
             �?������?�            �w@       x       �                    �?����[�?�            pp@       y       �                    �?�S����?z            �g@       z       �                    @L@\��1��?l            �d@       {       �                    �?���.�6�?X            @a@       |       �                   @E@Hn�.P��?N             _@        }       ~                    ]@      �?             @        ������������������������       �                     �?               �                   �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@(;L]n�?J             ^@        ������������������������       �                     �I@        �       �                   c@p��%���?*            @Q@        ������������������������       �                      @        �       �                   �b@0�,���?)            �P@       �       �                    �?0�z��?�?%             O@       ������������������������       �                     H@        �       �                   0k@@4և���?             ,@        �       �                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?d}h���?
             ,@       ������������������������       �                     "@        �       �                   �e@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �\@����X�?             <@        ������������������������       �                      @        �       �                    @M@�θ�?             :@        ������������������������       �                     @        �       �                   ps@�LQ�1	�?             7@       �       �                   0q@�C��2(�?             6@       �       �                    q@؇���X�?             ,@       �       �                    �M@$�q-�?
             *@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?r�q��?             8@       �       �                     Q@d}h���?	             ,@       �       �                   `^@�8��8��?             (@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     $@        �       �                     R@��pBI�?.            @R@       �       �                   s@�k~X��?-             R@       ������������������������       �        $             N@        �       �                    �?�8��8��?	             (@       ������������������������       �                     "@        �       �                   (s@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?���dQ'�?K            �\@        �       �                    �?؇���X�?            �A@       ������������������������       �                     9@        �       �                   �^@      �?             $@        �       �                   �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          `ff�?�o;����?6            �S@       �       �                    �?ؓ��M{�?!            �K@       �       �                   pb@D^��#��?            �D@        �       �                   �n@���!pc�?	             &@       �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �       	          @33�?      �?             @        ������������������������       �                      @        �       �                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?d��0u��?             >@        �       �                   �m@�C��2(�?             &@        ������������������������       �                     @        �       �                   0e@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�\��N��?             3@        ������������������������       �                     @        �       �                   a@�q�q�?	             .@       �       �                   �X@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �o@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?	             ,@       ������������������������       �                     (@        ������������������������       �                      @        �       �                   �`@r�q��?             8@        �       �                   �a@�z�G��?	             $@        ������������������������       �                     @        �       �                    �?և���X�?             @       �       �                   `d@�q�q�?             @       �       �                    �?�q�q�?             @       �       �       	             @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    ]@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �t�b�4     h�h*h-K ��h/��R�(KK�KK��ha�B0        u@     �x@     �G@     `o@      3@      5@      &@      @       @      @      �?              �?      @      �?       @               @      �?                      @      "@               @      0@      @      0@      @      �?              �?      @                      .@      @              <@     �l@      2@      S@      *@     �R@      @      *@      @      @              @      @      �?              �?      @                      "@       @      O@              2@       @      F@       @      >@              $@       @      4@      �?       @              @      �?      @               @      �?       @      �?                       @      @      (@               @      @      @      @               @      @              @       @      �?       @                      �?              ,@      @      �?      @              �?      �?      �?                      �?      $@     @c@      @     �P@      @      0@       @      0@      �?      0@              &@      �?      @      �?      �?      �?                      �?              @      �?               @              @     �I@       @              �?     �I@      �?      @              @      �?                      H@      @     �U@       @      T@      �?      T@      �?      .@      �?       @               @      �?                      *@             @P@      �?              �?      @              @      �?             r@     `b@      2@     �D@       @      6@      �?              �?      6@      �?      .@              (@      �?      @      �?                      @              @      0@      3@      0@      ,@      0@      @      (@       @      @              @       @               @      @              @      @       @      @              @       @      �?       @                      �?       @                       @              @     �p@     �Z@     �l@      @@      d@      >@     �b@      1@      `@      "@     �]@      @       @       @      �?              �?       @               @      �?              ]@      @     �I@             @P@      @               @     @P@       @     �N@      �?      H@              *@      �?       @      �?       @                      �?      &@              @      �?              �?      @              &@      @      "@               @      @              @       @              4@       @               @      4@      @              @      4@      @      4@       @      (@       @      (@      �?      �?      �?      �?                      �?      &@                      �?       @                      �?      &@      *@      &@      @      &@      �?      �?      �?      �?                      �?      $@                       @              $@     �Q@       @     �Q@      �?      N@              &@      �?      "@               @      �?              �?       @                      �?      D@     �R@      @      >@              9@      @      @      @      �?              �?      @               @      @      �?      @      �?                      @      �?             �A@      F@      ?@      8@      3@      6@       @      @       @      �?      @              @      �?       @              �?      �?      �?                      �?               @      &@      3@      �?      $@              @      �?      @              @      �?              $@      "@              @      $@      @       @       @              �?       @      �?      @              �?      �?      �?                      �?       @      @       @                      @      (@       @      (@                       @      @      4@      @      @              @      @      @       @      @       @      �?      �?      �?      �?                      �?      �?                      @      �?              �?      *@      �?                      *@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ	�tlhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B@-         P                    �?�+	G�?�           ��@                      
             �?�@o-4�?�            �s@                                 �g@P���Q�?y             i@                                 �O@��:x�ٳ?x            �h@      �?������������������������       �                     @                                  �a@`�E���?u            @h@      �?������������������������       �        %             O@                                  �a@Pa�	�?P            �`@        	       
                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �? g�yB�?N             `@                                  �?�x�E~�?8            @V@        ������������������������       �                    �E@                                  �e@�nkK�?             G@                                 @[@      �?             @@                                  @Y@      �?              @ �s��  ������������������������       �                     �?given RV������������������������       �                     �? y_like
                           �?(;L]n�?             >@y_like
                          �e@���7�?             6@see doc������������������������       �                     3@ ation)
                            H@�q�q�?             @ aramete������������������������       �                      @      s������������������������       �                     �? --
    ������������������������       �                      @on evalu������������������������       �                     ,@ r   r�������������������������       �                     D@ r   �������������������������       �                      @r�   r�       G                    �?�>4ևF�?G             \@  s"         *                    @K@�c�Α�?8            �U@                )                    �?l��[B��?             =@}tt!       &                    �?r�q��?             2@      @"       %                    �D@����X�?             @       #       $                    �?      �?             @      �?������������������������       �                      @        ������������������������       �                      @      @������������������������       �                     @      @'       (                     F@�C��2(�?
             &@       @������������������������       �                     �?      �?������������������������       �        	             $@      �?������������������������       �                     &@      �?+       D                    �?д>��C�?#             M@      @,       3                   pk@���@��?            �B@        -       .                    �?@4և���?
             ,@      �?������������������������       �                     "@      >@/       2       
             �?z�G�z�?             @     �?0       1                   �b@      �?             @       ������������������������       �                     @      8@������������������������       �                     �?        ������������������������       �                     �?        4       5                   �k@8����?             7@      $@������������������������       �                      @        6       ?       	          `ff�?���N8�?             5@       @7       >       
             �?���Q��?             @     �?8       =                    �?      �?             @       9       :                   @[@�q�q�?             @       @������������������������       �                     �?      @;       <                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        @       A                    �N@      �?             0@       ������������������������       �                     &@        B       C                   �`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        E       F                   `c@�����?             5@       ������������������������       �        
             3@        ������������������������       �                      @        H       O                    c@�+e�X�?             9@       I       J                   0n@�q�q�?             8@        ������������������������       �                     *@        K       L                    �?�eP*L��?             &@        ������������������������       �                     @        M       N                   �a@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        Q       �                    @.�����?           `z@       R       y       
             �?��4:���?�            Px@        S       t                     P@�a7���?4            �U@       T       U                   `X@x�(�3��?/            @S@        ������������������������       �                     @        V       q                    �?����>�?.            �R@       W       l                    �?     8�?&             P@       X       _                    �?��[�p�?            �G@        Y       Z                    �J@��
ц��?             *@        ������������������������       �                     @        [       ^                    �?      �?              @        \       ]                   �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        `       k                    @N@�t����?             A@       a       j                   �b@�C��2(�?            �@@       b       i                   @^@      �?             @@        c       h       	          @33�?�r����?	             .@       d       g                     E@@4և���?             ,@        e       f                   �h@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �                     �?        m       n                    @M@�IєX�?	             1@       ������������������������       �                     "@        o       p                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        r       s                   `\@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        u       v                    �?�����H�?             "@       ������������������������       �                     @        w       x                    `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        z       �                   �e@�č����?�            �r@       {       |       	          ����?�Tޫvɼ?�            �r@        ������������������������       �        !             L@        }       �                    �?� �$m�?�            �n@       ~                          �m@�����?�            �h@       ������������������������       �        D            �Z@        �       �                   �m@�ܸb���?<             W@        ������������������������       �                     @        �       �                    �R@����!p�?;             V@       �       �                    @M@`��F:u�?:            �U@       �       �                   �_@ �Jj�G�?$            �K@        �       �                   �\@@4և���?
             ,@        �       �                   �[@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                    �D@        �       �                    �M@     ��?             @@        �       �                   �`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �^@h�����?             <@        �       �                   �`@�8��8��?	             (@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        
             0@        ������������������������       �                     �?        �       �       	          ����?�3Ea�$�?"             G@        ������������������������       �                     @        �       �                    �Q@���H��?             E@       �       �       
             �?������?            �D@       �       �                   pc@������?             B@       ������������������������       �                    �@@        �       �                    �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   @^@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   pb@�eP*L��?            �@@       �       �                    �?X�<ݚ�?             ;@       �       �                    �?ҳ�wY;�?             1@       �       �                    �?8�Z$���?             *@       �       �                    �O@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �n@���Q��?             $@       �       �                   @`@      �?              @        �       �                   �i@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�BP       `t@     �y@      m@     �S@     �g@      $@     �g@       @              @     �g@      @      O@              `@      @      �?       @               @      �?             �_@       @     �U@       @     �E@              F@       @      >@       @      �?      �?      �?                      �?      =@      �?      5@      �?      3@               @      �?       @                      �?       @              ,@              D@                       @     �E@     @Q@      8@     �O@      ,@      .@      @      .@       @      @       @       @       @                       @              @      �?      $@      �?                      $@      &@              $@      H@       @      =@      �?      *@              "@      �?      @      �?      @              @      �?                      �?      @      0@       @              @      0@      @       @       @       @      �?       @              �?      �?      �?      �?                      �?      �?              �?               @      ,@              &@       @      @       @                      @       @      3@              3@       @              3@      @      3@      @      *@              @      @      @              �?      @              @      �?                      �?     @W@     �t@     �R@     �s@     �K@      ?@      K@      7@              @      K@      4@     �J@      &@     �B@      $@      @      @              @      @      �?       @      �?       @                      �?      @              >@      @      >@      @      >@       @      *@       @      *@      �?       @      �?              �?       @              &@                      �?      1@                      �?              �?      0@      �?      "@              @      �?              �?      @              �?      "@              "@      �?              �?       @              @      �?      �?              �?      �?              4@     �q@      2@     �q@              L@      2@     `l@      "@     �g@             �Z@      "@     �T@      @              @     �T@      @     �T@      �?      K@      �?      *@      �?      @              @      �?                      "@             �D@      @      =@       @       @               @       @              �?      ;@      �?      &@      �?      �?              �?      �?                      $@              0@      �?              "@     �B@      @              @     �B@      @     �B@      �?     �A@             �@@      �?       @               @      �?              @       @      @                       @      �?               @              2@      .@      (@      .@      @      &@       @      &@       @      "@              "@       @                       @      @              @      @      @       @      �?       @               @      �?              @                       @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�ޡhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKㅔh��B�8         `                    �?6������?�           ��@      &@       3       	          ����?v���a�?�            @r@               &                   �b@03�Z*!�?L            �^@      @                           �?� ���?@            @Z@      @                          �s@,sI�v�?8            �V@     �?              
             �?�Zl�i��?4            @T@      @                           �?�q�q�?             (@      @������������������������       �                     @        	       
       	          ����?�<ݚ�?             "@      �?������������������������       �                      @     �?������������������������       �                     @     &@                           \@�nkK�?-            @Q@      �?                          �k@�����?             5@     $@������������������������       �        
             0@                                   @K@���Q��?             @      �?������������������������       �                      @                                    P@�q�q�?             @     @������������������������       �                      @      @������������������������       �                     �?                      	          `ff�?@��8��?             H@      �?������������������������       �                     4@      7@                           @G@h�����?             <@      $@                           �?�����H�?             "@     �?������������������������       �                     @      @                          �`@�q�q�?             @      �?������������������������       �                      @        ������������������������       �                     �?      �?������������������������       �                     3@      �?                           �?�q�q�?             "@        ������������������������       �                     @      �?������������������������       �                     @      L@        !                   �\@��S���?             .@     �T@������������������������       �                     @      K@"       %                   `c@���!pc�?             &@       #       $                   @a@�����H�?             "@      @������������������������       �                      @      &@������������������������       �                     �?      $@������������������������       �                      @        '       2       	          ����?�q�q�?             2@    �@@(       1                    �?      �?
             0@      @)       0                    �?���Q��?             $@       *       +                    �?X�<ݚ�?             "@      &@������������������������       �                      @       @,       -                   @`@և���X�?             @       @������������������������       �                      @       @.       /                     M@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        4       ]                    @$�q-�?r             e@       5       6                   �U@��M6�?o            `d@        ������������������������       �                      @        7       <                    �?��	l�?n             d@        8       9                   �`@�<ݚ�?             "@        ������������������������       �                     @        :       ;                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        =       V                    �?@+K&:~�?h             c@       >       ?                   `]@��S�ۿ?>            �V@        ������������������������       �        	             ,@        @       U                    �R@�˹�m��?5             S@       A       T                    @N@��S�ۿ?4            �R@       B       M                    @M@h�WH��?&             K@       C       F                    �?�nkK�?!             G@        D       E       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        G       H                    �? qP��B�?            �E@       ������������������������       �                    �B@        I       J                   @_@r�q��?             @        ������������������������       �                     @        K       L                    �I@      �?              @  ��&� ������������������������       �                     �?        ������������������������       �                     �?        N       S                    o@      �?              @       O       P                   P`@r�q��?             @        ������������������������       �                     @        Q       R       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                     �?        W       \                    �?0�z��?�?*             O@       X       [                     K@����?�?            �F@        Y       Z                    ]@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@        ������������������������       �                     1@        ^       _                   �i@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        a       �                    �?�C�"��?"           �{@       b       �                    �?�1��u�?�            �v@       c       ~                    �?     ��?�             p@       d       q                    @L@Ά^���?e            �b@       e       j       
             �?�8��8��?P             ^@       f       g                    �? f^8���?D            �Y@       ������������������������       �        :            @V@        h       i                   `e@d}h���?
             ,@       ������������������������       �        	             &@        ������������������������       �                     @        k       n                    �F@j���� �?             1@        l       m       	             @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        o       p       
             �?���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        r       }                    �P@*;L]n�?             >@       s       z                    �?r�q��?             8@       t       y                    �O@���Q��?
             .@       u       x                   �`@      �?	             (@       v       w                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        {       |       	          ����?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               �                   pe@�ǧ\�?D            �Z@        �       �       
             �?���Q��?             9@       �       �                   @E@@4և���?             ,@        �       �                   @_@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                    `@"pc�
�?             &@        �       �                   @\@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�w���?5            @T@        �       �                    �?�P�*�?             ?@       �       �                    @L@����X�?             5@       �       �                    �D@@�0�!��?             1@        �       �                   �e@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @I@$�q-�?	             *@       ������������������������       �                     "@        �       �                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �f@�z�G��?             $@       �       �       	          @33�?      �?              @       �       �                   �[@r�q��?             @       �       �                   g@�q�q�?             @        ������������������������       �                     �?        �       �                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   c@�J�4�?             I@       �       �                    `@Pa�	�?            �@@       �       �                   �_@      �?             0@        ������������������������       �                      @        �       �                   @a@      �?              @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             1@        �       �                   �_@j���� �?	             1@       �       �                   �\@      �?              @        ������������������������       �                     @        �       �                    �H@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             "@       �       �                   �c@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `X@�~i��?G            @[@        �       �       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?�����?E            @Z@       �       �                   @c@pY���D�?2            �S@       ������������������������       �        .            �Q@        �       �                    �N@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �D@�	j*D�?             :@        ������������������������       �                      @        �       �       	          `ff@      �?             8@       ������������������������       �                     1@        �       �                    b@؇���X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?�w�r��?2            @S@        �       �                   �U@����e��?            �@@        ������������������������       �                     *@        ������������������������       �                     4@        �       �                   �k@��2(&�?             F@       �       �                    �?XB���?             =@       ������������������������       �                     9@        �       �                    b@      �?             @       �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   pm@�q�q�?	             .@        ������������������������       �                     @        �       �       	          ����?�C��2(�?             &@       ������������������������       �                     "@        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B0       �t@     �x@      F@      o@      ?@      W@      3@     �U@      &@     �S@       @     @R@      @      @      @               @      @       @                      @      @     �P@       @      3@              0@       @      @               @       @      �?       @                      �?      �?     �G@              4@      �?      ;@      �?       @              @      �?       @               @      �?                      3@      @      @      @                      @       @      @              @       @      @       @      �?       @                      �?               @      (@      @      (@      @      @      @      @      @       @              @      @               @      @       @      @                       @      �?              @                       @      *@     �c@      &@      c@       @              "@      c@       @      @              @       @      @              @       @              @      b@      @      U@              ,@      @     �Q@      @     �Q@      @     �H@       @      F@      �?       @      �?                       @      �?      E@             �B@      �?      @              @      �?      �?              �?      �?              @      @      �?      @              @      �?       @      �?                       @       @                      5@      �?              �?     �N@      �?      F@      �?      @      �?                      @              C@              1@       @      @       @                      @     0r@     �b@     �p@      Y@      e@      V@     �_@      7@     �[@      $@      Y@      @     @V@              &@      @      &@                      @      $@      @      @      �?      @                      �?      @      @              @      @              1@      *@      &@      *@      "@      @      "@      @      @      @              @      @              @                      @       @      @       @                      @      @             �D@     @P@      .@      $@      *@      �?      @      �?      �?      �?              �?      �?               @              $@               @      "@       @       @               @       @                      @      :@     �K@      2@      *@      .@      @      ,@      @       @       @       @                       @      (@      �?      "@              @      �?      @                      �?      �?      @              @      �?              @      @      �?      @      �?      @      �?       @              �?      �?      �?              �?      �?                      @               @       @               @      E@      �?      @@      �?      .@               @      �?      @      �?      �?              �?      �?                      @              1@      @      $@      �?      @              @      �?      @              @      �?              @      @      @      �?      @               @      �?       @                      �?               @     @X@      (@       @       @       @                       @     �W@      $@     @S@       @     �Q@              @       @               @      @              2@       @               @      2@      @      1@              �?      @              �?      �?      @      �?                      @      :@     �I@      4@      *@              *@      4@              @      C@      �?      <@              9@      �?      @      �?      �?              �?      �?                       @      @      $@      @              �?      $@              "@      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJQY%hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKՅ�h��B@5         f                    �?�Z���?�           ��@                                   �?$��n�?�             s@ 0,N,0,U              	          433�?      �?             0@    �P@              
             �?ףp=
�?             $@      @������������������������       �                     "@        ������������������������       �                     �?                                  �`@r�q��?             @     �?������������������������       �                     @        	       
                     K@�q�q�?             @ |f|j������������������������       �                     �?�|f������������������������       �                      @dd| j       O                    �?���7��?�             r@|� |              
             �?�iX/�1�?�            �n@ D �\|                           c@8^s]e�?             =@dd�|                          �g@������?             ;@ | jd
d������������������������       �                     "@k�rN|                          pq@b�2�tk�?             2@      @                           �?��
ц��?             *@     �B@������������������������       �                     @      �?                          �i@�q�q�?             "@      @������������������������       �                      @                                   �?؇���X�?             @     F@������������������������       �                     @      C@������������������������       �                     �?      @������������������������       �                     @      7@������������������������       �                      @      @       N                    �R@��ҘR�?�             k@     �?       5                   pa@���Hx�?�             k@     @                          �h@ d���W�?s            @f@      @������������������������       �        /            �Q@               4                    �?88��M�?D            �Z@               !                   pi@����1�?2            @R@      $@������������������������       �                     �?      �?"       +       	          ����?�8��8��?1             R@      "@#       $                    @K@�<ݚ�?             2@      @������������������������       �                     &@      @%       &                   �`@և���X�?             @      �?������������������������       �                     @      �?'       *                    �?      �?             @     @(       )                    @M@      �?              @      �?������������������������       �                     �?      @������������������������       �                     �?      @@������������������������       �                      @      �?,       -       	          ���@ 7���B�?%             K@     1@������������������������       �                     F@      @.       /                   8p@z�G�z�?             $@      �?������������������������       �                     @      �?0       3                    `@�q�q�?             @        1       2       	          ���@�q�q�?             @        ������������������������       �                      @       @������������������������       �                     �?      @������������������������       �                     @      @������������������������       �                     A@        6       M                    �?p�ݯ��?             C@     @7       F                   �n@|��?���?             ;@      @8       9       	          @33�?�����?             3@      "@������������������������       �                     �?        :       E                   �b@�E��ӭ�?             2@       ;       <                    U@X�Cc�?	             ,@        ������������������������       �                     @        =       D                   �\@      �?             $@       >       C       	          ��� @����X�?             @       ?       @                    �?���Q��?             @        ������������������������       �                     �?        A       B                   �m@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        G       H                   �p@      �?              @        ������������������������       �                     @        I       L                    �?      �?             @       J       K                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        P       _                   �`@�eP*L��?             F@        Q       ^                    �?�z�G��?
             4@       R       S                   �Z@�<ݚ�?	             2@        ������������������������       �                     �?        T       W                   �j@@�0�!��?             1@        U       V                    `@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        X       Y                    �?�C��2(�?             &@        ������������������������       �                     @        Z       [                    @I@r�q��?             @        ������������������������       �                     @        \       ]                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        `       a       
             �?      �?             8@        ������������������������       �                     @        b       e                    �H@ףp=
�?             4@        c       d       	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             0@        g       �       	          pff�?~�Q7:�?           �z@       h       �       
             �?x�X9���?�            �u@       i       j       	          033�     ��?�             p@        ������������������������       �                     @        k       �                    �?$%j����?�            �o@       l                          �g@�1��?o            �e@       m       |                    �?��+��<�?n            �e@       n       w       	            �?���tcH�?L            @^@       o       p                    @G@�ջ����?C             Z@        ������������������������       �        !             J@        q       r                   n@ pƵHP�?"             J@       ������������������������       �                     @@        s       v                    �H@P���Q�?             4@        t       u                   @c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        x       {                   @b@������?	             1@        y       z                   @a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        }       ~                     R@���J��?"            �I@       ������������������������       �        !             I@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @D@R���Q�?0             T@        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��G���?,            �R@       �       �                   @E@      �?#             L@        �       �                    �?���Q��?             @        �       �                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �c@�:�]��?            �I@       ������������������������       �                     B@        �       �                   �i@������?             .@        ������������������������       �                     @        �       �       	          `ff�?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �?b�2�tk�?	             2@       �       �                    q@���|���?             &@        �       �                   8p@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?
��^���?9            @W@        �       �                    c@���Q��?             >@       �       �                   �\@ �o_��?             9@        ������������������������       �                     @        �       �                    �?"pc�
�?             6@       �       �       	          ����?�	j*D�?	             *@       �       �       	          ����?      �?              @       �       �       	          ����?�q�q�?             @       �       �                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �       	          hff�?�[|x��?&            �O@       ������������������������       �                     H@        �       �                     P@�q�q�?	             .@       �       �                    \@      �?             $@        ������������������������       �                     @        �       �                   �W@����X�?             @        �       �                   �s@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��qC�?9            �S@       �       �                    �?д>��C�?+             M@        �       �       	             �?�	j*D�?             :@        ������������������������       �                     �?        �       �                   pb@ �o_��?             9@       �       �                   �o@�GN�z�?             6@       �       �                   �a@�q�q�?             .@        ������������������������       �                     @        �       �                   m@X�<ݚ�?             "@       �       �                    �N@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@      �?             @@       ������������������������       �                     :@        �       �                     M@�q�q�?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���N8�?             5@        ������������������������       �                     &@        �       �                    b@      �?             $@        ������������������������       �                     @        �       �                    @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�BP        u@     �x@     �N@     �n@      $@      @      "@      �?      "@                      �?      �?      @              @      �?       @      �?                       @     �I@     �m@      ?@     �j@      "@      4@      @      4@              "@      @      &@      @      @      @              @      @       @              �?      @              @      �?                      @       @              6@     `h@      5@     `h@      @     `e@             �Q@      @      Y@      @     �P@      �?              @     �P@      @      ,@              &@      @      @      @              �?      @      �?      �?      �?                      �?               @       @      J@              F@       @       @              @       @      @       @      �?       @                      �?              @              A@      ,@      8@      ,@      *@      *@      @              �?      *@      @      "@      @      @              @      @      @       @      @       @              �?      @      �?      @                      �?       @                      @      @              �?      @              @      �?      @      �?      �?              �?      �?                       @              &@      �?              4@      8@      ,@      @      ,@      @              �?      ,@      @      @       @               @      @              $@      �?      @              @      �?      @              �?      �?      �?                      �?               @      @      2@      @               @      2@       @       @       @                       @              0@     Pq@     �b@     `o@     �X@     �l@      <@              @     �l@      9@     �d@      @     �d@      @      ]@      @     �Y@      �?      J@             �I@      �?      @@              3@      �?      @      �?              �?      @              ,@              *@      @      @      @      @                      @      "@              I@      �?      I@                      �?              �?      O@      2@       @      @              @       @              N@      ,@     �H@      @       @      @      �?      �?      �?                      �?      �?       @               @      �?             �G@      @      B@              &@      @              @      &@      �?      &@                      �?      &@      @      @      @      @      @              @      @                      @      @              7@     �Q@      2@      (@      2@      @              @      2@      @      "@      @      @      @      @       @      �?       @      �?                       @      @                       @      @              "@                      @      @      M@              H@      @      $@      @      @              @      @       @      �?       @               @      �?              @                      @      :@     �J@      $@      H@       @      2@      �?              @      2@      @      1@      @      $@              @      @      @       @      @              @       @              @                      @       @      �?              �?       @               @      >@              :@       @      @       @      �?       @                      �?              @      0@      @      &@              @      @      @               @      @              @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��fbhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B@/         R                    �?�#i����?�           ��@      �?              
             �?�� ~E��?�            s@0,Up,0       
                    I@�8��8��?y            �i@     �m@                           ^@8�Z$���?             *@      "@������������������������       �                     �?                                 Pb@�8��8��?             (@     �?������������������������       �                     "@               	                    �J@�q�q�?             @      �?������������������������       �                      @        ������������������������       �                     �?                                   @L@�w��3(�?s            �g@                                 @[@���=��?]            �b@                                   �?�C��2(�?             &@        ������������������������       �                     @                                  �Z@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        X            `a@      �?              	          833@,���i�?            �D@     1@                          p@$�q-�?            �C@      @������������������������       �                     7@      &@                          �c@     ��?	             0@    �p@                          @a@�q�q�?             "@       ������������������������       �                     @      Z@������������������������       �                     @      I@������������������������       �                     @      @������������������������       �                      @      =@       /                    �?:�o���?@            @Y@               (                   �a@������?            �F@              '                    �?PN��T'�?             ;@     @                           �k@�<ݚ�?             2@        ������������������������       �                     "@      @!       &                   �b@X�<ݚ�?             "@       "       #       	             �?r�q��?             @     �?������������������������       �                     @       @$       %       	             �?�q�q�?             @      @������������������������       �                     �?      �?������������������������       �                      @      @������������������������       �                     @     �Q@������������������������       �                     "@      @)       .       	          ����?X�<ݚ�?             2@       @*       -                    �N@���!pc�?             &@      @+       ,                   @_@z�G�z�?             $@      M@������������������������       �                      @      @������������������������       �                      @        ������������������������       �                     �?      H@������������������������       �                     @      1@0       M       	          ��� @      �?&             L@     @1       J                   �b@~���L0�?            �H@     @2       C                    �?���N8�?             E@     >@3       B                    �?�û��|�?             7@       4       5                    @F@�\��N��?             3@        ������������������������       �                     @      @6       ;                   �l@�	j*D�?
             *@        7       8                   @_@      �?              @       ������������������������       �                     @        9       :                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        <       A       
             �?���Q��?             @       =       @                    �?      �?             @       >       ?                   @_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        D       E                   �`@�}�+r��?             3@       ������������������������       �                     (@        F       I                   �`@؇���X�?             @        G       H                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     @        K       L                   �^@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        N       O       	          `ff@؇���X�?             @        ������������������������       �                     @        P       Q                   @L@      �?             @        ������������������������       �                     �?       ������������������������       �                     @        S       �       
             �?�f|��?           �z@        T       ]                    P@H�౅z�?R            �`@        U       V                    [@r�q��?             >@        ������������������������       �                     �?        W       \                    �?\-��p�?             =@        X       [                    a@և���X�?             @        Y       Z                   @^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        ^       }       	          ����?�ެD��?A            �Y@       _       l                    �L@��܂O�?8            �V@       `       g                   @\@85�}C�?#            �N@        a       f                    �F@������?             .@       b       c                   �i@���Q��?             $@        ������������������������       �                      @        d       e                    �E@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @       h       i                   �b@��<b�ƥ?             G@       ������������������������       �                     E@        j       k                   po@      �?             @        ������������������������       �                     �?       ������������������������       �                     @       m       n                    �?*;L]n�?             >@        ������������������������       �                     @       o       v                    �?�q�q�?             8@       p       q                   �b@r�q��?             2@       ������������������������       �                     &@       r       u                    @և���X�?             @       s       t                   @d@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        w       |                   f@�q�q�?             @       x       y                   0a@z�G�z�?             @        ������������������������       �                     @       z       {                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?       ~       �                    �?      �?	             (@              �                   �d@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @K@����8�?�            �r@        �       �                    �? ��+,��?P            @_@       �       �       
             �?�h����?G             \@       �       �                    �?`�߻�ɒ?C             [@       ������������������������       �        2            �T@        �       �                    �G@`2U0*��?             9@        �       �                   �i@z�G�z�?             @       ������������������������       �                     @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    @H@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �H@8�Z$���?	             *@       �       �                     E@�q�q�?             @        ������������������������       �                     @        �       �                   �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �a@��Sa+��?x            `e@        �       �       	          033�?p���?"             I@       ������������������������       �                     =@        �       �                    �?���N8�?             5@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             1@        �       �       
             �?"pc�
�?V            @^@       �       �                   Pi@�՘���?F            �W@        �       �                    �?���!pc�?             &@       �       �                   `]@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?r�q��??             U@        �       �                    �?և���X�?             <@       �       �                   pm@�eP*L��?             6@        ������������������������       �                     @        �       �                   �^@�q�q�?             .@        �       �                    _@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                   Xw@h�����?,             L@       �       �                    �O@@3����?*             K@       ������������������������       �                    �C@        �       �                   �a@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        �       �                   0c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �t�b��      h�h*h-K ��h/��R�(KK�KK��ha�B�       `u@     �x@     @m@     �Q@     `g@      1@       @      &@      �?              �?      &@              "@      �?       @               @      �?              g@      @     �b@      �?      $@      �?      @              @      �?      @                      �?     `a@              B@      @      B@      @      7@              *@      @      @      @      @                      @      @                       @     �G@      K@      (@     �@@      @      7@      @      ,@              "@      @      @      �?      @              @      �?       @      �?                       @      @                      "@       @      $@       @      @       @       @               @       @                      �?              @     �A@      5@      A@      .@      @@      $@      ,@      "@      $@      "@      @              @      "@      �?      @              @      �?      �?      �?                      �?      @       @       @       @      �?       @               @      �?              �?              �?              @              2@      �?      (@              @      �?      �?      �?      �?                      �?      @               @      @       @                      @      �?      @              @      �?      @      �?                      @      [@     t@     @T@      J@      @      9@      �?              @      9@      @      @      �?      @      �?                      @      @                      6@      S@      ;@     @R@      2@      L@      @      &@      @      @      @               @      @       @      @                       @      @             �F@      �?      E@              @      �?              �?      @              1@      *@              @      1@      @      .@      @      &@              @      @      �?      @              @      �?              @               @      @      �?      @              @      �?      �?      �?                      �?      �?              @      "@      �?      "@              "@      �?               @              ;@     �p@      @     @^@       @     �[@      �?     �Z@             �T@      �?      8@      �?      @              @      �?      �?      �?                      �?              4@      �?      @              @      �?               @      &@       @      @              @       @      �?              �?       @                      @      7@     �b@      �?     �H@              =@      �?      4@      �?      @              @      �?                      1@      6@     �X@      6@     @R@       @      @      @      �?              �?      @              �?       @               @      �?              ,@     �Q@      (@      0@      (@      $@      @              @      $@      @      �?              �?      @                      "@              @       @      K@      �?     �J@             �C@      �?      ,@              ,@      �?              �?      �?              �?      �?                      :@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ$�phG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKÅ�h��B�0         P       
             �?"��G,�?�           ��@      &@       A                    �?DE��2{�?�            �r@p,0
39                           �?6C�d�?�            �o@     �?              	             @Pq�����?m            @e@                                 �g@�|�%T�?l             e@                                  �?h�����?k             e@     @              	            �? �h�7W�?C            �Z@     @                          @[@`Ӹ����?9            �V@      @	       
                   �Z@�q�q�?             "@      @������������������������       �                     @      "@������������������������       �                     @       @                          �t@ �)���?5            @T@     5@������������������������       �        4             T@      "@������������������������       �                     �?      @                          @a@      �?
             0@       @������������������������       �                      @                                  @b@      �?              @        ������������������������       �                      @      @������������������������       �                     @        ������������������������       �        (             O@      8@������������������������       �                     �?      @������������������������       �                     �?      �?       *                   �j@��]�T��?2            �T@      �?       '                    i@�eP*L��?            �@@     2@       &                    �?�q�q�?             8@                                  �?�G��l��?             5@    �X@                           @L@ףp=
�?             $@     @������������������������       �                     @                                   �M@�q�q�?             @      �?������������������������       �                     �?      @������������������������       �                      @                !                    �H@"pc�
�?             &@      �?������������������������       �                     @     @^@"       #                   @Z@���Q��?             @      8@������������������������       �                      @        $       %                     P@�q�q�?             @     @������������������������       �                      @      @������������������������       �                     �?      @������������������������       �                     @      4@(       )                    _@�����H�?             "@      1@������������������������       �                     �?      �?������������������������       �                      @       @+       <                   �b@ \� ���?            �H@     $@,       /                    �?�T|n�q�?            �E@      �?-       .                    �?���Q��?             @     K@������������������������       �                     @      ,@������������������������       �                      @        0       3                   `\@�KM�]�?             C@        1       2                   p`@      �?             @        ������������������������       �                     @        ������������������������       �                     @        4       ;       	          ����?      �?             @@       5       6                    �?P���Q�?             4@       ������������������������       �                     $@        7       :                   f@ףp=
�?             $@       8       9                    �L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        =       >                   Hq@r�q��?             @        ������������������������       �                     @        ?       @                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        B       O       	          `ff�?r�q��?             H@       C       D                    �?¦	^_�?             ?@        ������������������������       �        	             .@        E       F                   @V@     ��?
             0@        ������������������������       �                     @        G       L       	          833�?��
ц��?	             *@        H       K                    �H@r�q��?             @        I       J                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        M       N                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             1@        Q       j                   �g@�*�@P��?            {@        R       c                   0b@�Km�a̾?T            �a@       S       `                   �c@X�?٥�??            �Y@       T       U                    �?`�(c�?;            �X@       ������������������������       �        #             M@        V       _                    �?��(\���?             D@        W       Z                    �J@r�q��?             2@        X       Y       
             �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        [       \                   Pb@$�q-�?             *@       ������������������������       �                     $@        ]       ^                    �P@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@       a       b                   0d@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @       d       i                    �P@������?            �B@       e       f                    �? >�֕�?            �A@       ������������������������       �                     >@        g       h                    �?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        k       t                    �?d}h���?�            `r@        l       m                   Pl@r�q��?             8@        ������������������������       �                     @       n       s                    b@ҳ�wY;�?
             1@       o       p                   �p@      �?             (@        ������������������������       �                     @        q       r                    �?؇���X�?             @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @        u       �                    @�+$�jP�?�            �p@       v       �                   �a@>��k�	�?�            �o@       w       �                    �?��o�x,�?a            �c@       x       �                    �?6kh�h��?T            �`@       y       �                    �?�Y�?�(�?A            �[@       z       �                    m@h��Q(�?%            �P@        {       |                    @K@�5��?             ;@        ������������������������       �                     (@        }       �       
             �?������?             .@       ~                           �L@d}h���?             ,@        ������������������������       �                      @        �       �                    `@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    _@��(\���?             D@        ������������������������       �                     7@        �       �                    `@@�0�!��?             1@        ������������������������       �                      @        �       �                    @M@��S�ۿ?             .@       ������������������������       �        	             *@        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �J@�Ra����?             F@        �       �       	              @      �?              @       �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @M@������?             B@        �       �                    c@��S�ۿ?             .@       ������������������������       �        	             *@        �       �                    [@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �       �                   �Z@�û��|�?             7@        ������������������������       �                     @        �       �                    �?�z�G��?             4@        �       �                    ]@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?r�q��?
             (@        �       �                    `@      �?             @        ������������������������       �                     �?        �       �                   �u@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���}<S�?             7@       ������������������������       �                     ,@        �       �       
             �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?p�qG�?4             X@        �       �                   �_@�חF�P�?             ?@       ������������������������       �        	             *@        �       �                   @b@�E��ӭ�?             2@        ������������������������       �                     @        �       �                   `c@�q�q�?             (@        �       �       	             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        #            @P@        �       �                    �?j���� �?
             1@       �       �                   0`@�q�q�?             "@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     P@      �?              @        ������������������������       �                     @        �       �                    �P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B0       @s@     �z@     �m@      P@     �j@      C@     @d@       @     @d@      @     @d@      @      Y@      @     �U@      @      @      @      @                      @      T@      �?      T@                      �?      ,@       @       @              @       @               @      @              O@                      �?              �?      J@      >@      .@      2@      ,@      $@      &@      $@      "@      �?      @               @      �?              �?       @               @      "@              @       @      @               @       @      �?       @                      �?      @              �?       @      �?                       @     �B@      (@      B@      @       @      @              @       @              A@      @      @      @      @                      @      ?@      �?      3@      �?      $@              "@      �?      @      �?      @                      �?      @              (@              �?      @              @      �?      �?      �?                      �?      6@      :@      6@      "@      .@              @      "@              @      @      @      �?      @      �?       @      �?                       @              @      @      �?              �?      @                      1@      R@     �v@      "@     ``@      @     �X@      @     �W@              M@      @     �B@      @      .@       @      @              @       @              �?      (@              $@      �?       @               @      �?                      6@       @      @       @                      @      @     �@@       @     �@@              >@       @      @       @                      @       @             �O@     �l@      *@      &@      @              @      &@      @      @              @      @      �?              �?      @                      @      I@     �k@      D@     �j@     �A@     �^@     �@@     @Y@      3@      W@      ,@     �J@      &@      0@              (@      &@      @      &@      @       @              @      @              @      @                      �?      @     �B@              7@      @      ,@       @              �?      ,@              *@      �?      �?      �?                      �?      @     �C@      @      @      �?      @              @      �?              @              �?     �A@      �?      ,@              *@      �?      �?      �?                      �?              5@      ,@      "@              @      ,@      @      @      @       @               @      @              @       @              $@       @       @       @              �?       @      �?       @                      �?       @               @      5@              ,@       @      @              @       @              @     �V@      @      :@              *@      @      *@              @      @      @      @      �?              �?      @                      @             @P@      $@      @      @      @      @      �?      @                      �?              @      @      �?      @               @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJW:+LhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKم�h��B@6         N                   �`@�#i����?�           ��@       @                           �?p�L���?�            `s@ M,NAP,1              
             �?����X�?             <@     �?������������������������       �                     4@        ������������������������       �                      @       @       #       
             �?&Eȧ��?�            �q@       @              	          ����?�ݏ^���?             �F@                                   �?z�G�z�?             4@     �?	                           @�<ݚ�?             2@      @
                          �]@     ��?
             0@      "@������������������������       �                     $@       @                           W@      �?             @      5@������������������������       �                     @      "@������������������������       �                     @      @                           ^@      �?              @       @������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @      @                           �? �o_��?             9@      @������������������������       �                     @      1@                           �?"pc�
�?             6@    �W@                           _@�C��2(�?	             &@     @������������������������       �                     "@      $@                          �_@      �?              @      6@������������������������       �                     �?     �@@������������������������       �                     �?                       	          033�?���!pc�?             &@     &@                          @\@؇���X�?             @      @������������������������       �                     @      @                           �?      �?              @     @Y@������������������������       �                     �?      (@������������������������       �                     �?      @!       "                    S@      �?             @     �B@������������������������       �                      @      ,@������������������������       �                      @      �?$       ?                    �?\ ���?�            �m@     @%       &                   i@P�9�׸?u             f@      ,@������������������������       �        -            �N@      �?'       (                   @i@ج��w�?H            �\@      @������������������������       �                     �?      @)       >                    �?l�b�G��?G            �\@     �?*       7       	          ����?�^;\��?5            @V@        +       6                   `^@R�}e�.�?             :@     @,       -                    `@     ��?             0@      *@������������������������       �                     @      �?.       5                   �]@�	j*D�?	             *@    @P@/       0                    @K@"pc�
�?             &@        ������������������������       �                     @        1       4                    �L@�q�q�?             @       2       3                    b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        8       =                   �_@ ������?%            �O@        9       <                   pp@ףp=
�?             $@       :       ;                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �J@        ������������������������       �                     9@        @       A                   �k@L=�m��?'            �N@       ������������������������       �                     B@        B       M       	             @� �	��?             9@       C       D                   �_@���|���?             6@        ������������������������       �                      @        E       L                   `c@և���X�?             ,@       F       G                     N@�eP*L��?             &@        ������������������������       �                     @        H       I                    �O@؇���X�?             @        ������������������������       �                     @        J       K       	          @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        O       �       
             �?������?
           �z@       P       �       	          ���@d��cό�?�             o@       Q       f                    �?����B��?�            �n@       R       Y                   @[@�d���?l            �e@        S       T                     F@r�q��?             @        ������������������������       �                     @       U       X                    �?�q�q�?             @       V       W                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     �?        Z       e                   �c@�h����?f             e@        [       b                   �c@Ћ����?1            �T@       \       a                    _@�Fǌ��?/            �S@        ]       ^                   (p@h�����?             <@       ������������������������       �                     8@        _       `                   �^@      �?             @       ������������������������       �                     @       ������������������������       �                     �?        ������������������������       �                     �I@        c       d                     M@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @       ������������������������       �        5            �U@        g       �                    �?��
P�?-            �Q@       h       }       	          hff�?��H�}�?              I@       i       n                    f@�E��ӭ�?             B@        j       m                    �?      �?              @       k       l                   Pe@      �?             @       ������������������������       �                     @        ������������������������       �                     @       ������������������������       �                      @       o       x                    �L@�>4և��?             <@       p       w       	          ����?�8��8��?             8@       q       r                    �I@ףp=
�?             4@       ������������������������       �                     *@       s       t                   Pc@����X�?             @        ������������������������       �                     @        u       v                    @K@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?       ������������������������       �                     @       y       z                   p`@      �?             @        ������������������������       �                      @        {       |                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ~       �                    @և���X�?	             ,@              �                    b@���!pc�?             &@       �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �M@P���Q�?             4@       ������������������������       �        
             1@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�tp��\�?m            �e@       �       �                    �?      �?Y             b@       �       �                   �r@�^�X�?:            @X@       �       �                   o@�E��ӭ�?6            �V@       �       �       	          `ff�?�5��?#             K@       �       �                    �?�4�����?             ?@        ������������������������       �                     @        �       �       	          ����?���Q��?             9@        ������������������������       �                     @        �       �                    @�X����?             6@       �       �                   �g@p�ݯ��?             3@        �       �                   `c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @d@d}h���?	             ,@       �       �                    @E@r�q��?             (@        ������������������������       �                     �?        �       �                    b@�C��2(�?             &@        �       �       	          ����?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�nkK�?             7@       ������������������������       �                     2@        �       �                   @^@z�G�z�?             @        ������������������������       �                      @        �       �       	             @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�8��8��?             B@        �       �                    �I@      �?             (@       ������������������������       �                      @        �       �                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     8@        �       �                   @_@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?z�J��?            �G@        �       �                   �q@r�q��?             8@       �       �                   �g@P���Q�?             4@        �       �                    �?�q�q�?             @       �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             1@        �       �                   �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �a@�㙢�c�?             7@        �       �                    �?���Q��?             $@       �       �                    �?      �?              @       �       �                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@        �       �                    �?��� ��?             ?@        ������������������������       �        	             *@        �       �       	          `ff@�<ݚ�?             2@       �       �       
             �?      �?
             0@       �       �                   �c@r�q��?             (@       ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       `u@     �x@     �O@     �n@      4@       @      4@                       @     �E@     �m@      7@      6@      0@      @      ,@      @      *@      @      $@              @      @              @      @              �?      �?      �?                      �?       @              @      2@      @              @      2@      �?      $@              "@      �?      �?      �?                      �?      @       @      �?      @              @      �?      �?              �?      �?               @       @       @                       @      4@      k@      "@     �d@             �N@      "@     �Z@      �?               @     �Z@       @     @T@      @      3@      @      "@      @              @      "@       @      "@              @       @      @       @      �?       @                      �?              @       @                      $@      �?      O@      �?      "@      �?      @              @      �?                      @             �J@              9@      &@      I@              B@      &@      ,@       @      ,@               @       @      @      @      @      @              �?      @              @      �?       @      �?                       @      @              @             pq@      b@     �k@      <@     �k@      7@     @e@      @      @      �?      @               @      �?      �?      �?              �?      �?              �?             �d@      @     �S@      @     �S@      �?      ;@      �?      8@              @      �?      @                      �?     �I@              �?       @      �?                       @     �U@             �I@      3@      @@      2@      :@      $@      @      @      @      @      @                      @               @      7@      @      6@       @      2@       @      *@              @       @      @              �?       @               @      �?              @              �?      @               @      �?      �?              �?      �?              @       @      @       @      �?       @              @      �?       @      �?                       @       @              @              3@      �?      1@               @      �?       @                      �?              @      M@     @]@      K@     �V@      >@     �P@      9@     @P@      6@      @@      5@      $@      @              .@      $@              @      .@      @      (@      @      �?      @              @      �?              &@      @      $@       @              �?      $@      �?      @      �?      @                      �?      @              �?      �?      �?                      �?      @              �?      6@              2@      �?      @               @      �?       @      �?                       @      @     �@@      @      "@               @      @      �?      @                      �?              8@      @       @      @                       @      8@      7@      4@      @      3@      �?       @      �?      �?      �?      �?                      �?      �?              1@              �?      @      �?                      @      @      3@      @      @       @      @      �?      @      �?                      @      �?       @               @      �?               @                      *@      @      ;@              *@      @      ,@       @      ,@       @      $@              @       @      @       @                      @              @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJF<KdhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKǅ�h��B�1         X       
             �?�#i����?�           ��@                                   U@4>���?�             u@        ������������������������       �                     @      @       '                    �?����s��?�            �t@                                  I@��ɶ�"�?�            �i@       @       	                    �Q@     ��?             0@     @                          �d@r�q��?             (@     d@������������������������       �                     $@      N@������������������������       �                      @        
                           �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @               &                    �?�F�l���?y            �g@                                 @[@ >�֕�?W            �a@                                  `m@���|���?             &@        ������������������������       �                     @                                   @I@և���X�?             @        ������������������������       �                     @      @������������������������       �                     @      @                          pa@0Ƭ!sĮ?Q             `@     1@                           �?@�z�G�?4             T@    �W@                           �?@3����?#             K@      @                          p@ �q�q�?             8@     $@������������������������       �                     4@      6@                          �_@      �?             @     �@@                          Pr@      �?              @        ������������������������       �                     �?     &@������������������������       �                     �?      @������������������������       �                      @      @������������������������       �                     >@     @Y@������������������������       �                     :@      (@        %                   �a@��<D�m�?            �H@     @!       "                    �N@ܷ��?��?             =@      @������������������������       �                     9@        #       $                   @t@      �?             @      @������������������������       �                     �?     @P@������������������������       �                     @      $@������������������������       �                     4@      @������������������������       �        "            �I@       @(       O                    �?     x�?L             `@       )       D                   �b@Rg��J��?;            �X@       *       9       	          ����?0�� ��?(            �O@     2@+       4                   @E@�KM�]�?             C@        ,       -                    �?      �?             @       @������������������������       �                      @      8@.       /                    �?      �?             @      7@������������������������       �                     �?      �?0       1                   `Y@�q�q�?             @        ������������������������       �                     �?      3@2       3                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?      *@5       8                   `_@      �?             @@      @6       7                    @r�q��?             @     @������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@        :       ;                   @^@���Q��?             9@        ������������������������       �                     @        <       C                    �?      �?             4@       =       >       	          ����?�q�q�?	             (@        ������������������������       �                     @        ?       @                     N@����X�?             @        ������������������������       �                     @        A       B                   0k@�q�q�?             @       ������������������������       �                      @       ������������������������       �                     �?        ������������������������       �                      @        E       N                    f@4�2%ޑ�?            �A@       F       M       	          ����?"pc�
�?            �@@       G       H                   ``@�����?             3@        ������������������������       �                     @        I       L                    @      �?             (@       J       K                     M@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                      @       P       W                    @�r����?             >@       Q       R                   �U@"pc�
�?             6@        ������������������������       �                      @        S       T                    s@ףp=
�?             4@       ������������������������       �                     ,@       U       V                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @       Y       �                    �?L�~m��?           �x@       Z       e                   �a@hh<>�?�            �q@        [       d                    �?��p\�?            �D@        \       a                   p`@�θ�?             *@       ]       `                    @K@      �?              @        ^       _                   �Z@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?       ������������������������       �                     @        b       c                    �L@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @       ������������������������       �                     <@       f       �       	          pff�?������?�             n@        g       �                    @lG:<�?<            @X@       h                          �a@\Ќ=��?9            �V@       i       v                    �? {��e�?             �J@       j       u                    �?��(\���?             D@       k       l       	          ����?ȵHPS!�?             :@        ������������������������       �                     ,@        m       n                    @K@      �?             (@        ������������������������       �                     @       o       p                   �[@      �?             @        ������������������������       �                      @       q       r       	          `ff�?      �?             @        ������������������������       �                      @       s       t                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@       w       ~                    �?�n_Y�K�?             *@       x       y                   p@���!pc�?             &@        ������������������������       �                     @        z       }                    �L@      �?             @       {       |       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �                      @       ������������������������       �                      @       �       �       	          ����?P����?             C@       �       �                    �D@������?             >@        ������������������������       �                     @        �       �                    �?8�Z$���?             :@        ������������������������       �                     @        �       �                   �m@�㙢�c�?             7@       �       �                   @_@���|���?             &@        �       �                    �F@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	            �?���Q��?             @       �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        �       �                   @`@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@r�q��?             @        ������������������������       �                     @        �       �                   `c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��K˱F�?c            �a@       �       �                   �b@L�'�7��?O            @]@       �       �                   �\@@uvI��?C            �X@        �       �                    �K@�C��2(�?             &@       ������������������������       �                     @        �       �       	             @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        >            �U@        �       �                    �?�\��N��?             3@        ������������������������       �                      @        �       �       	             @j���� �?
             1@       �       �                    e@����X�?             ,@       �       �                   0c@ףp=
�?             $@        �       �                   c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �e@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��
ц��?             :@        �       �                    �?ףp=
�?             $@        �       �       	          pff�?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     P@     ��?             0@       ������������������������       �        
             *@        ������������������������       �                     @        �       �                   �h@��x$�?G            �\@        ������������������������       �        "            �J@        �       �       	          ����?Hn�.P��?%             O@       �       �       	          ����?l��\��?             A@        ������������������������       �                     &@        �       �                    �P@�LQ�1	�?             7@       �       �                   i@�C��2(�?             6@        ������������������������       �                     �?        �       �                    �M@���N8�?             5@       ������������������������       �                     0@        �       �       	          ����?z�G�z�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     <@        �t�bh�h*h-K ��h/��R�(KK�KK��ha�Bp       `u@     �x@      q@     �P@              @      q@     �O@     @h@      *@      &@      @      $@       @      $@                       @      �?      @      �?                      @     �f@       @     �`@       @      @      @      @              @      @              @      @             @_@      @     �S@      �?     �J@      �?      7@      �?      4@              @      �?      �?      �?              �?      �?               @              >@              :@              G@      @      :@      @      9@              �?      @      �?                      @      4@             �I@             �S@      I@      J@      G@      F@      3@      A@      @      @      @       @              �?      @              �?      �?       @              �?      �?      �?      �?                      �?      ?@      �?      @      �?      @                      �?      :@              $@      .@      @              @      .@      @      @              @      @       @      @              �?       @               @      �?                       @       @      ;@      @      ;@      @      *@              @      @      @      @      @      @                      @              @              ,@       @              :@      @      2@      @               @      2@       @      ,@              @       @      @                       @       @             �Q@     `t@     �P@     �j@      @      C@      @      $@      �?      @      �?       @               @      �?                      @       @      @              @       @                      <@      P@      f@     �D@      L@      B@     �K@      &@      E@      @     �B@      @      7@              ,@      @      "@              @      @      @       @              �?      @               @      �?      �?      �?                      �?              ,@       @      @       @      @      @              @      @      �?      @              @      �?               @                       @      9@      *@      6@       @              @      6@      @      @              3@      @      @      @      @      �?      @                      �?       @      @       @      �?              �?       @                       @      (@              @      @      @                      @      @      �?      @               @      �?              �?       @              7@      ^@      &@     �Z@      �?     @X@      �?      $@              @      �?      @      �?                      @             �U@      $@      "@               @      $@      @      $@      @      "@      �?      �?      �?      �?                      �?       @              �?      @              @      �?                      @      (@      ,@      "@      �?      @      �?              �?      @              @              @      *@              *@      @              @      \@             �J@      @     �M@      @      ?@              &@      @      4@       @      4@      �?              �?      4@              0@      �?      @      �?       @      �?                       @               @      �?                      <@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJؽ�hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKŅ�h��B@1         H                    �?�/�$�y�?�           ��@     �U@              
             �?�V��Q�?�            0s@,ATA,14       
                    @L@��.N"Ҭ?|            �i@     @       	                    �? J���#�?f             f@                                 h@�K}��?<            �Y@     �?������������������������       �        :            �X@                                   d@      �?             @        ������������������������       �                     @      .@������������������������       �                     �?      k@������������������������       �        *            �R@                      	          @33�?�חF�P�?             ?@     "@                           �?ܷ��?��?             =@     @                          �s@@�0�!��?             1@     �?                           �?      �?             0@     O@                           �?r�q��?	             (@                                 @a@ףp=
�?             $@     I@������������������������       �                     @       @              	          @33�?�q�q�?             @      @������������������������       �                     �?       @                           �?      �?              @      <@������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?              @      �?������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @      2@������������������������       �                     �?        ������������������������       �                     (@       @������������������������       �                      @               )                   �`@
�c�Z�?B             Y@               &                    �?`�H�/��?            �I@     �?        %                   P`@��S�ۿ?            �F@       @!       "                   �\@؇���X�?             5@       ������������������������       �                     0@        #       $                    �?���Q��?             @     �?������������������������       �                     @      @������������������������       �                      @        ������������������������       �                     8@      ^@'       (                    �P@�q�q�?             @     @������������������������       �                     @     �U@������������������������       �                      @      @*       E       	             @�`���?%            �H@     �?+       2                    �I@H�z�G�?             D@        ,       /                    �?j���� �?             1@      �?-       .                   �\@����X�?             @      *@������������������������       �                      @     �J@������������������������       �                     @      4@0       1                     F@z�G�z�?             $@      0@������������������������       �                      @       @������������������������       �                      @        3       D                    �P@8����?             7@       4       5                   @J@���N8�?             5@        ������������������������       �                     �?        6       ?       	          ����?z�G�z�?             4@        7       >                    �?և���X�?             @       8       =       
             �?      �?             @       9       :                   l@���Q��?             @        ������������������������       �                     �?        ;       <                    ]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        @       A                   @m@$�q-�?
             *@        ������������������������       �                      @        B       C                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @       ������������������������       �                      @       F       G       
             �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?       I       |       	          ����?GI2�J�?           �z@        J       o                    �?���Q��?c             b@       K       f       
             �?Ć��H��?K            �Z@       L       a                    �?�j�'�=�?-            �P@       M       Z                    �?�&!��?!            �E@       N       Q                    �?V�a�� �?             =@        O       P                    b@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        R       W       	          ����?�C��2(�?             6@       S       V                    @D@�}�+r��?             3@        T       U                    a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        X       Y                    V@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        [       `                    �L@d}h���?
             ,@       \       ]                   g@և���X�?             @        ������������������������       �                      @        ^       _                   �p@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        b       c                    �?���}<S�?             7@       ������������������������       �                     1@        d       e                    s@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        g       h       	          833�?�p ��?            �D@       ������������������������       �                     ?@        i       j                   �X@���Q��?             $@        ������������������������       �                      @        k       l                    �?      �?              @        ������������������������       �                     �?        m       n                    @I@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        p       y                   �`@�?�'�@�?             C@       q       x                    �? �q�q�?             8@        r       s                   �^@�����H�?             "@       ������������������������       �                     @        t       u                   @a@�q�q�?             @        ������������������������       �                     �?        v       w                   �t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        z       {                   ``@����X�?	             ,@       ������������������������       �                     $@        ������������������������       �                     @        }       �                    �R@Tri����?�            �q@       ~       �                   h@ �Cc}�?�            �q@               �                   P`@�x�E~�?8            @V@       ������������������������       �        *             Q@        �       �       
             �?�����?             5@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@        �       �                   0i@�m	{�?u            �g@        �       �                    @�<ݚ�?             "@        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @ȵHPS!�?q            �f@       �       �                    _@�� ND��?h            `e@        �       �                   �\@�<ݚ�?             B@        �       �                    �J@�q�q�?             (@        �       �       	             @r�q��?             @       �       �                    Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?      �?             8@        ������������������������       �                     @        �       �                    @G@r�q��?             2@       �       �                    �?և���X�?             @       �       �                   `a@�q�q�?             @        ������������������������       �                     @        �       �                   �Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �       
             �?���?T            �`@        �       �                   �`@�E��ӭ�?             2@        ������������������������       �                     @        �       �                   �a@�q�q�?	             (@        �       �       	          ��� @      �?             @       �       �       	          033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@      �?              @        ������������������������       �                     @        �       �                   0l@      �?             @        ������������������������       �                     �?        �       �                    b@�q�q�?             @       �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �Q@ ���J��?H            @]@        ������������������������       �                     �?        �       �       	          ����? _�@�Y�?G             ]@        �       �                    �?�����?             5@       ������������������������       �                     *@        �       �                    �?      �?              @       �       �                    @O@�q�q�?             @       �       �                    @K@�q�q�?             @        ������������������������       �                     �?        �       �                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        9            �W@        �       �                    �?�eP*L��?	             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�b�M	     h�h*h-K ��h/��R�(KK�KK��ha�BP        t@     �y@     �l@     @S@      i@      @     �e@      �?     @Y@      �?     �X@              @      �?      @                      �?     �R@              :@      @      :@      @      ,@      @      ,@       @      $@       @      "@      �?      @               @      �?      �?              �?      �?              �?      �?              �?      �?      �?                      �?      @                      �?      (@                       @      =@     �Q@      @      G@      @      E@      @      2@              0@      @       @      @                       @              8@       @      @              @       @              8@      9@      7@      1@      @      $@      @       @               @      @               @       @       @                       @      0@      @      0@      @              �?      0@      @      @      @      @      @       @      @      �?              �?      @      �?                      @      �?              �?              (@      �?       @              @      �?              �?      @                       @      �?       @               @      �?             �V@     u@      M@     �U@     �J@      K@     �G@      3@      :@      1@      7@      @      @      @              @      @              4@       @      2@      �?       @      �?       @                      �?      0@               @      �?              �?       @              @      &@      @      @               @      @       @      @                       @              @      5@       @      1@              @       @      @                       @      @     �A@              ?@      @      @               @      @       @              �?      @      �?              �?      @              @     �@@      �?      7@      �?       @              @      �?       @              �?      �?      �?      �?                      �?              .@      @      $@              $@      @              @@     @o@      >@     @o@       @     �U@              Q@       @      3@       @      �?       @                      �?              2@      <@     `d@      @       @      �?       @      �?                       @      @              5@      d@      0@     `c@       @      <@      @      @      @      �?       @      �?              �?       @              @                      @      @      5@              @      @      .@      @      @       @      @              @       @      �?              �?       @              �?                      &@       @     �_@      @      *@              @      @      @      @      �?      �?      �?      �?                      �?       @               @      @              @       @       @              �?       @      �?      �?      �?      �?                      �?      �?              @     �\@      �?               @     �\@       @      3@              *@       @      @       @      @       @      �?      �?              �?      �?      �?                      �?              @               @             �W@      @      @              @      @               @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJX��vhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKŅ�h��B@1         X       
             �?���
%�?�           ��@                                   �?�˱��H�?�            �r@      @                          �j@
j*D>�?             J@      @                           �M@H%u��?             9@      �?������������������������       �                     ,@     �?       	                   �]@���!pc�?             &@                                   @N@      �?             @        ������������������������       �                      @      .@������������������������       �                      @      �?
                           �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @      �?                           �B@l��
I��?             ;@      �?������������������������       �                      @      @                           �L@�+e�X�?             9@     @                          d@�����H�?	             2@     �?������������������������       �                     &@                                  @d@����X�?             @        ������������������������       �                      @      3@������������������������       �                     @      @                          �p@և���X�?             @     �?              	          433�?���Q��?             @      �?������������������������       �                     @      @������������������������       �                      @       @������������������������       �                      @       @                          @V@��k�c��?�            `o@      ?@������������������������       �                      @      �?       7                    �?�5U��K�?�             o@    �@@       4                     R@Hx�i�.�?{             g@      @       )                    �? �ղ?y            �f@     �?       &                   h@ �Jj�G�?D            �[@               %                    _@`�߻�ɒ?B             [@      Q@!       $                    �?����?�?            �F@     �?"       #                   �^@��Y��]�?            �D@      @������������������������       �                     D@      d@������������������������       �                     �?      �?������������������������       �                     @        ������������������������       �        (            �O@      .@'       (                    d@      �?              @      �?������������������������       �                     �?      &@������������������������       �                     �?      @*       3       	          hff@���;QU�?5            @R@     �?+       0                    �O@0z�(>��?3            �Q@      @,       /                   @[@Pa�	�?/            �P@        -       .                    �?�q�q�?             @        ������������������������       �                      @      @������������������������       �                     @      �?������������������������       �        ,             N@       @1       2                   0b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        5       6                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        8       O       	          ����?      �?)             P@       9       H                    q@���B���?!             J@       :       =                    T@�L���?            �B@        ;       <                    [@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        >       E                    �?�IєX�?             A@       ?       @                   �e@h�����?             <@       ������������������������       �                     9@        A       D                    @�q�q�?             @       B       C                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        F       G                    @F@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        I       J                   �_@��S���?             .@        ������������������������       �                     @        K       N                    �?�����H�?             "@       L       M                    �I@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        P       W                    �?      �?             (@        Q       R                    k@؇���X�?             @        ������������������������       �                     @        S       T                    �?      �?             @        ������������������������       �                      @        U       V                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Y       �                    �? ��7E��?           �z@       Z       �                   �b@�����?�            `v@       [       \                   �U@�<� w�?�            �s@        ������������������������       �                     �?        ]       h                    �F@�u���?�            �s@        ^       _                   pf@"pc�
�?             6@        ������������������������       �                     "@        `       a                   �a@�	j*D�?	             *@        ������������������������       �                     @        b       g                    �?X�<ݚ�?             "@       c       f                    o@r�q��?             @        d       e                    �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        i       �       
             �?��P�/a�?�            pr@       j       w                    �?�Ń��̧?�            �o@        k       l                    @M@Hn�.P��?#             O@        ������������������������       �                     @@        m       v       	          ����?ףp=
�?             >@        n       u                   `@�θ�?	             *@       o       t                    �?�C��2(�?             &@       p       q                   �q@r�q��?             @       ������������������������       �                     @        r       s                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             1@        x       �       	          ����?���̅ӟ?|            �g@        y       z                   0l@ ��WV�?1            �S@       ������������������������       �                    �I@        {       �                   �`@�����H�?             ;@       |       }                   �l@�8��8��?             8@        ������������������������       �                     �?        ~       �       	          ����?�nkK�?             7@               �       	          ����?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        	             *@        �       �                    �?�q�q�?             @       �       �                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        K             \@        �       �                   �r@X�EQ]N�?            �E@       �       �                    �?��p\�?            �D@       ������������������������       �                     A@        �       �                    �?և���X�?             @        �       �       	             @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	          033�?�G�z�?             D@        �       �       
             �?      �?             0@       ������������������������       �        	             *@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             8@       �       �                    �?      �?
             0@        �       �                    �L@      �?              @       ������������������������       �                     @        �       �                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	             @      �?              @       �       �                   @_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     K@      �?              @        ������������������������       �                     @        �       �                     O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�!�,�E�?+            @R@        �       �                    �J@��a�n`�?             ?@        �       �                    �?���|���?             &@       �       �                   h@X�<ݚ�?             "@        ������������������������       �                      @        �       �                   �s@և���X�?             @       �       �                   `a@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             4@        �       �       	          ���@և���X�?             E@       �       �                    �?�t����?             A@       �       �                    �?؇���X�?             <@       �       �                    c@P���Q�?             4@        ������������������������       �                     &@        �       �                   �b@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �F@      �?              @        ������������������������       �                      @        �       �                   0l@r�q��?             @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�BP       0s@     �z@     �n@      L@      6@      >@      @      6@              ,@      @       @       @       @       @                       @      �?      @      �?                      @      3@       @               @      3@      @      0@       @      &@              @       @               @      @              @      @      @       @      @                       @               @      l@      :@               @      l@      8@      f@       @      f@      @      [@       @     �Z@      �?      F@      �?      D@      �?      D@                      �?      @             �O@              �?      �?      �?                      �?      Q@      @      Q@      @      P@       @      @       @               @      @              N@              @      �?      @                      �?               @      �?      �?      �?                      �?      H@      0@      E@      $@      A@      @       @      �?       @                      �?      @@       @      ;@      �?      9@               @      �?      �?      �?              �?      �?              �?              @      �?              �?      @               @      @              @       @      �?      @      �?      @                      �?      @              @      @      �?      @              @      �?      @               @      �?      �?      �?                      �?      @              N@     0w@      =@     �t@      0@     �r@      �?              .@     �r@      @      2@              "@      @      "@              @      @      @      �?      @      �?      �?              �?      �?                      @      @              &@     �q@      @     �n@      @     �M@              @@      @      ;@      @      $@      �?      $@      �?      @              @      �?      �?      �?                      �?              @       @                      1@      @     `g@      @     �R@             �I@      @      8@       @      6@      �?              �?      6@      �?      "@              "@      �?                      *@      �?       @      �?      �?              �?      �?                      �?              \@      @      C@      @      C@              A@      @      @      @      �?      @                      �?              @       @              *@      ;@      �?      .@              *@      �?       @      �?                       @      (@      (@      $@      @      @      �?      @               @      �?       @                      �?      @      @      @      �?              �?      @                      @       @      @              @       @      �?       @                      �?      ?@      E@      @      8@      @      @      @      @       @              @      @      �?      @              @      �?               @               @                      4@      8@      2@      8@      $@      8@      @      3@      �?      &@               @      �?       @                      �?      @      @               @      @      �?       @      �?       @                      �?      @                      @               @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���EhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKǅ�h��B�1         R       	          033�?�r,��?�           ��@     6@       /       
             �?H;N	�	�?�             x@                                 @E@8Ӈ���?�            `p@      @                          @^@8�A�0��?             6@       @������������������������       �                     @     �G@                          `V@���Q��?             .@      @������������������������       �                      @      3@       	                    �J@��
ц��?
             *@      @������������������������       �                     @      @
                          �]@      �?              @      "@������������������������       �                     @       @                          `_@���Q��?             @      5@������������������������       �                      @      "@������������������������       �                     @      @                           �?��(\���?�             n@      @                          �t@��8����?}             h@                                 d@�~��?y            �f@       ������������������������       �        L             \@                                  Pd@����Q8�?-            �Q@      �?                          0o@      �?             @     @������������������������       �                     @       @������������������������       �                     @                                  �b@ ����?)            @P@       ������������������������       �        %            �M@      "@                           �?r�q��?             @     �?������������������������       �                     @        ������������������������       �                     �?      @@                          u@�����H�?             "@      @������������������������       �                     �?      �?������������������������       �                      @     `g@       (                    q@r�qG�?              H@     6@        %                     P@�t����?             A@     "@!       "                    �? 7���B�?             ;@     �?������������������������       �                     5@      \@#       $                   �j@r�q��?             @      @������������������������       �                     �?      @������������������������       �                     @      *@&       '                    �P@և���X�?             @      (@������������������������       �                     @      �?������������������������       �                     @      �?)       .       	          @33�?X�Cc�?
             ,@     @*       -                   (s@      �?             (@     �?+       ,                    �?ףp=
�?             $@      @������������������������       �                     �?      @������������������������       �                     "@      4@������������������������       �                      @      �?������������������������       �                      @      �?0       5                   �g@�&�5y�?J             _@      �?1       4                    �?`���i��?             F@      @2       3                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �D@        6       =                   �a@��Q��?.             T@        7       8                   0i@l��\��?             A@        ������������������������       �                     �?        9       :       	          ����?�FVQ&�?            �@@       ������������������������       �                     :@        ;       <                   �m@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        >       C                   @^@�LQ�1	�?             G@        ?       B                    �?�q�q�?             .@       @       A                    �?�θ�?             *@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        D       Q                    �?�n`���?             ?@       E       P                    �?\-��p�?             =@       F       G       	          ����?������?	             1@        ������������������������       �                      @        H       O       
             �?�r����?             .@       I       J                    �J@؇���X�?             ,@        ������������������������       �                     �?        K       N                    �L@$�q-�?             *@        L       M                   Pj@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        S       �                   P`@д>��C�?�            �u@        T       �                    �?�w�"w��?e             c@       U       V                    V@�n`���??            @W@        ������������������������       �                     �?        W       �                   �b@��H�?>             W@       X              
             �?�p ��?9            �T@       Y       j                    @L@�Y����?0            �P@       Z       i                   �_@��-�=��?            �C@       [       \                   �h@\-��p�?             =@        ������������������������       �                     *@        ]       ^                   �Y@      �?             0@        ������������������������       �                     @        _       d                    �I@�	j*D�?
             *@        `       a                   �\@      �?             @        ������������������������       �                      @        b       c                   `]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        e       h                    �J@�����H�?             "@        f       g       	              @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        k       t                    ^@����X�?             <@        l       s                    �?X�<ݚ�?             "@       m       n                    �?և���X�?             @        ������������������������       �                     �?        o       r                   `]@      �?             @       p       q                   �X@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        u       ~                    @�S����?             3@       v       w       	          033�?�����H�?             2@        ������������������������       �                     @        x       y                   �_@"pc�
�?
             &@        ������������������������       �                     �?        z       }       
             �?ףp=
�?	             $@        {       |                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             .@        �       �                    �?      �?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@f�<�>��?&            �M@        �       �                    @O@�<ݚ�?             ;@       �       �                    �?�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?        �       �                    �O@X�<ݚ�?             "@        ������������������������       �                     @        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    W@     ��?             @@        ������������������������       �                     @        �       �       	          ����?�q�q�?             ;@       �       �       	          033�?D�n�3�?             3@       �       �                   �d@d}h���?
             ,@       �       �                   �b@ףp=
�?             $@        �       �       	          033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �p@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @B@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          pff�?�)���Y�?w            �h@       �       �                   �c@�חF�P�?=            @W@       �       �                    `@��(\���?3             T@       ������������������������       �        #            �J@        �       �                    �?�<ݚ�?             ;@        �       �                   ``@@4և���?             ,@        �       �                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                     P@�n_Y�K�?             *@       �       �                    �?X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�	j*D�?
             *@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                   �c@      �?             @       �       �                     F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?      �?             @        ������������������������       �                      @        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    `P@ f^8���?:            �Y@       �       �                   �a@��f�{��?/            �U@        �       �                   pa@�(\����?             D@        ������������������������       �        
             5@        �       �                    �?�}�+r��?
             3@       ������������������������       �                     1@        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     G@        �       �                    �?�t����?             1@       ������������������������       �        
             .@        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�Bp       �t@     Py@     �p@     @]@     `m@      ;@      *@      "@      @              @      "@               @      @      @              @      @       @      @              @       @               @      @             �k@      2@     `g@      @     `f@      @      \@             �P@      @      @      @              @      @              P@      �?     �M@              @      �?      @                      �?       @      �?              �?       @             �A@      *@      >@      @      :@      �?      5@              @      �?              �?      @              @      @              @      @              @      "@      @      "@      �?      "@      �?                      "@       @               @              A@     �V@      �?     �E@      �?       @               @      �?                     �D@     �@@     �G@      @      ?@      �?               @      ?@              :@       @      @       @                      @      >@      0@      @      $@      @      $@      @                      $@       @              9@      @      9@      @      *@      @               @      *@       @      (@       @              �?      (@      �?      @      �?      @                      �?       @              �?              (@                       @      N@      r@      E@     �[@      2@     �R@      �?              1@     �R@      (@     �Q@      (@     �K@      @     �A@      @      9@              *@      @      (@              @      @      "@      @      �?       @              �?      �?      �?                      �?      �?       @      �?       @               @      �?                      @              $@       @      4@      @      @      @      @              �?      @      @      �?      @      �?                      @       @               @              @      0@       @      0@              @       @      "@      �?              �?      "@      �?       @               @      �?                      @      �?                      .@      @      @      @                      @      8@     �A@      @      5@      �?      1@              1@      �?              @      @      @               @      @       @                      @      2@      ,@              @      2@      "@      &@       @      &@      @      "@      �?      �?      �?      �?                      �?       @               @       @               @       @                      @      @      �?              �?      @              2@     @f@      .@     �S@      @     �R@             �J@      @      5@      �?      *@      �?      @              @      �?                      $@      @       @      @      @      @                      @              @      "@      @      @              @      @      �?      @      �?       @      �?                       @              �?      @      �?       @              �?      �?              �?      �?              @      Y@      �?     @U@      �?     �C@              5@      �?      2@              1@      �?      �?      �?                      �?              G@       @      .@              .@       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ:9)bhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hK
hxK�hyh*h-K ��h/��R�(KK���h��B�.         N                    �?T8���?�           ��@      �?       7                    �?�s�ۺ�?�             s@                     	          ����?�3Ea�$�?n             g@       @              
             �?���Q��?            �F@      @                          �V@r�q��?             2@       @������������������������       �                     �?       @                           �?�t����?
             1@      @       	                    �?"pc�
�?             &@      @������������������������       �                     @    on a
                          @`@      �?             @ changed������������������������       �                     �?1.2.

                            �d@�q�q�?             @ eprecat������������������������       �                     �?ter : in������������������������       �                      @erform.
������������������������       �                     @e machin              	          ����?�����H�?             ;@    Cho������������������������       �                     7@      @                          �\@      �?             @       @������������������������       �                     �?      �?������������������������       �                     @               (                   P`@hb����?T            `a@     �[@       #                    �?P̏����?!            �L@    �Q@                          �U@�����H�?            �F@      *@������������������������       �                     �?      �?                           �b@�C��2(�?             F@     �?                           �M@�(\����?             D@       ������������������������       �                     :@      @                          `]@@4և���?             ,@      @������������������������       �                     @                                  �Z@؇���X�?             @      "@������������������������       �                     �?       @������������������������       �                     @      .@!       "       	             �?      �?             @     �A@������������������������       �                     �?        ������������������������       �                     @        $       %                   �n@      �?             (@      "@������������������������       �                     @      �?&       '       	          ����?      �?             @       @������������������������       �                     @      �?������������������������       �                     @     �S@)       6                    @������?3            �T@     *@*       +       	          `ff�? 7���B�?2            @T@     $@������������������������       �                    �H@      @,       1                   �a@     ��?             @@      @-       0                   k@      �?              @       @.       /                    �?�q�q�?             @      �?������������������������       �                     �?     @U@������������������������       �                      @      1@������������������������       �                     @      G@2       3       
             �? �q�q�?             8@       ������������������������       �                     6@        4       5                     Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        8       G                    �?�.�?�P�?Q             ^@       9       F                   hp@ '��h�?I            @[@       :       C                   @b@86��Z�?1            �S@       ;       >       
             �?��
���?-            �R@        <       =                    c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       B                    �G@`����֜?*            �Q@        @       A                    �F@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        &            �N@        D       E                   �a@      �?             @       ������������������������       �                     @       ������������������������       �                     �?        ������������������������       �                     >@        H       M                   �a@�eP*L��?             &@       I       L       	          ����?؇���X�?             @       J       K                   �_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        O       �       	          ����?�yZ����?           �z@       P       u       
             �?j�!����?�            0s@       Q       Z                   @E@���ܩm�?�            @m@        R       Y                    �?�eP*L��?             6@       S       T                    �?����X�?             ,@        ������������������������       �                     @       U       X                   @_@      �?              @       V       W       	          @33�?z�G�z�?             @        ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     @       ������������������������       �                      @       [       t                   �g@ T͋�x�?�            �j@       \       e                    �?��
�j�?�            @j@       ]       ^                    @L@��惡�?d             d@       ������������������������       �        R             `@        _       `                   �a@     ��?             @@        ������������������������       �        	             2@        a       b                   p@d}h���?	             ,@        ������������������������       �                      @        c       d                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     @        f       k                    �?ZՏ�m|�?            �H@       g       h                   �b@�7��?            �C@       ������������������������       �                     B@        i       j                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        l       q                   @_@���Q��?             $@       m       n                   �c@z�G�z�?             @        ������������������������       �                      @        o       p                   0l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        r       s                   �b@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @       v       w                   �`@X~�pX��?.            @R@        ������������������������       �                     3@        x       �                    �?���3L�?!             K@        y       �       
             �?z�G�z�?             4@       z       {                   @\@����X�?
             ,@        ������������������������       �                     �?        |                          �a@�θ�?	             *@        }       ~                    a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?              @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          833�?H�V�e��?             A@       �       �                    @h�����?             <@       ������������������������       �                     4@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?v�2t5�?Q            �^@       �       �                   �c@VP��g��?=             W@       �       �                   8w@�8��8��?(             N@       �       �       	          ����? ,��-�?'            �M@        �       �                   @Z@      �?             (@        ������������������������       �                     @   � � �       �                    �?      �?              @       �       �                   �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?`Ql�R�?            �G@        �       �                     G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �E@        ������������������������       �                     �?        �       �                    U@     ��?             @@        �       �                    �?����X�?             @       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?z�G�z�?             9@       �       �                    �L@�IєX�?             1@       ������������������������       �        	             *@        �       �                    @M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pe@      �?              @       �       �                    @z�G�z�?             @       �       �                   �d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @N@��a�n`�?             ?@       �       �                   `c@��S�ۿ?             .@       ������������������������       �        
             ,@        ������������������������       �                     �?        �       �       	          ���@      �?	             0@       �       �                   �]@r�q��?             (@        �       �                    `P@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       �t@     @y@     �G@     p@      B@     �b@      2@      ;@      .@      @              �?      .@       @      "@       @      @               @       @              �?       @      �?              �?       @              @              @      8@              7@      @      �?              �?      @              2@     @^@      ,@     �E@      @      D@      �?              @      D@      �?     �C@              :@      �?      *@              @      �?      @      �?                      @      @      �?              �?      @              "@      @      @              @      @      @                      @      @     �S@      @     �S@             �H@      @      =@       @      @       @      �?              �?       @                      @      �?      7@              6@      �?      �?              �?      �?              �?              &@     @[@      @      Z@      @     �R@       @     @R@      �?      @              @      �?              �?     @Q@      �?       @               @      �?                     �N@      @      �?      @                      �?              >@      @      @      @      �?      @      �?              �?      @               @                      @     �q@     `b@      m@     �R@      j@      9@      $@      (@      $@      @      @              @      @      �?      @      �?                      @      @                       @     �h@      *@     �h@      &@     �c@      @      `@              =@      @      2@              &@      @       @              @      @              @      @             �D@       @     �B@       @      B@              �?       @               @      �?              @      @      �?      @               @      �?       @               @      �?              @       @      @                       @               @      7@      I@              3@      7@      ?@      0@      @      $@      @              �?      $@      @      @       @      @                       @      @      �?      �?      �?      �?                      �?      @              @              @      ;@      �?      ;@              4@      �?      @              @      �?              @             �I@      R@      ;@     @P@      @     �K@      @     �K@      @      "@              @      @      @      @      �?              �?      @                      @      �?      G@      �?      @      �?                      @             �E@      �?              6@      $@       @      @              @       @       @               @       @              4@      @      0@      �?      *@              @      �?              �?      @              @      @      �?      @      �?      @      �?                      @              �?      @              8@      @      ,@      �?      ,@                      �?      $@      @      $@       @       @       @               @       @               @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�BHzhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKӅ�h��B�4         V       	          ����?�[��N�?�           ��@      ;@       1       
             �?��)��?�            �v@0,N,0,U                          `^@0�|#�p�?�            �o@      �?                           �?V������?            �B@     8@                           �?���}<S�?             7@      $@������������������������       �                     @                                   �?�����H�?             2@       ������������������������       �                      @      �?	       
                   �]@z�G�z�?             $@     �?������������������������       �                      @        ������������������������       �                      @                                   \@X�Cc�?             ,@     �V@������������������������       �                     @                                   @"pc�
�?             &@                                 �_@ףp=
�?             $@       ������������������������       �                     @      $@                           �?      �?             @      �?������������������������       �                     @      @������������������������       �                     �?        ������������������������       �                     �?     �R@       0                   h@��g�?~            @k@                     	          ���ٿp)�����?}             k@      @������������������������       �                      @      &@       /                    �?� Λ��?|            �j@              .       	            �?��'#��?X            �b@     @                           �?���D�k�?Q            �`@                                 @[@      �?:             X@      @������������������������       �                      @       @                          �t@��K2��?9            �W@      @������������������������       �        8            @W@      ?@������������������������       �                     �?      @        !                    T@���@��?            �B@      �?������������������������       �                      @        "       %                    �?b�h�d.�?            �A@      4@#       $                   `m@���Q��?             @        ������������������������       �                     @     �K@������������������������       �                      @      �?&       +                   �q@�r����?             >@     G@'       (                   @c@HP�s��?             9@    �E@������������������������       �        
             3@      @)       *                   �i@�q�q�?             @      @������������������������       �                      @      �?������������������������       �                     @      @,       -                   Pe@���Q��?             @       ������������������������       �                     @      �?������������������������       �                      @       @������������������������       �                     .@        ������������������������       �        $            �P@        ������������������������       �                      @        2       ?       	          ����?��>4��?H             \@       3       4                   Pi@(�s���?7             U@        ������������������������       �                    �@@        5       :                    �?`�H�/��?            �I@        6       7                   �n@և���X�?             @        ������������������������       �                     @        8       9                   �_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ;       <                    �?`���i��?             F@       ������������������������       �                    �A@        =       >                    @O@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        @       M                    �?      �?             <@       A       F                    �?      �?	             (@       B       C                   �\@؇���X�?             @       ������������������������       �                     @        D       E                     L@�q�q�?             @        ������������������������       �                     �?G D�&� ������������������������       �                      @        G       H                   Pa@���Q��?             @        ������������������������       �                     �?        I       L                    �?      �?             @       J       K                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        N       Q                    `@     ��?             0@        O       P       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        R       S                    �?�C��2(�?             &@       ������������������������       �                     @        T       U                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        W       �                    �?ByL5���?�            �v@       X       �                    �?���?�            ps@       Y       �                    @�W�a=�?�            �l@       Z       e       
             �?4�0_���?�            @l@        [       `                    S@�X����?             6@        \       ]                     M@և���X�?             @        ������������������������       �                      @        ^       _                   @_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        a       d                   �`@z�G�z�?             .@        b       c       	          `ff�?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        f       u       	          ����?�K��?|            �i@        g       r                   pb@�LQ�1	�?             G@       h       i                   �i@�7��?            �C@       ������������������������       �                     6@        j       k                    �?�t����?             1@        ������������������������       �                     "@        l       q                   �`@      �?              @       m       p                    �?؇���X�?             @       n       o                   �j@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        s       t                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        v       �                    _@�;u�,a�?`            �c@        w       x                    �H@������?            �B@        ������������������������       �                     (@        y       �                    �?�J�4�?             9@       z       �                    �?����X�?	             ,@       {       �       	          `ff�?r�q��?             (@        |       }                    �?      �?             @        ������������������������       �                     �?        ~                           @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        �       �                   �K@ ��+&ɐ?J            @^@        �       �       	          ����?�IєX�?             1@        �       �       	          033�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �        ?             Z@        �       �                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@�<ݚ�?8            @T@       �       �                     D@4և����?$             L@        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �Q@�NW���?"            �J@        �       �                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����? "��u�?              I@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?�nkK�?             G@       �       �                    �? ���J��?            �C@       ������������������������       �                     =@        �       �                    ^@ףp=
�?             $@        �       �                    �Q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @P@؇���X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    e@�q�����?             9@       �       �                   �^@������?             .@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	            �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    @C@z�G�z�?             $@        ������������������������       �                     �?        �       �       
             �?�����H�?             "@        �       �                    �?�q�q�?             @       �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �R@���>4��?(             L@        ������������������������       �                     @        �       �       
             �?�q�����?$             I@        ������������������������       �                     (@        �       �                    �?p�ݯ��?             C@       �       �                   h@�㙢�c�?             7@        ������������������������       �                      @        �       �                    _@�����?             5@        �       �                    Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�}�+r��?             3@        ������������������������       �                     $@        �       �                     N@�����H�?             "@       ������������������������       �                     @        �       �                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �n@�q�q�?             .@        �       �                   `c@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     P@և���X�?             @       �       �                   �x@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KK�KK��ha�B0       �s@     Pz@      o@     �]@     �l@      :@      :@      &@      5@       @      @              0@       @       @               @       @       @                       @      @      "@      @               @      "@      �?      "@              @      �?      @              @      �?              �?             `i@      .@     `i@      *@               @     `i@      &@      a@      &@     �^@      &@     @W@      @               @     @W@      �?     @W@                      �?      =@       @               @      =@      @      @       @      @                       @      :@      @      7@       @      3@              @       @               @      @              @       @      @                       @      .@             �P@                       @      3@     @W@      @     �S@             �@@      @      G@      @      @      @              �?      @              @      �?              �?     �E@             �A@      �?       @               @      �?              ,@      ,@      @      "@      �?      @              @      �?       @      �?                       @       @      @      �?              �?      @      �?      �?              �?      �?                       @      &@      @      �?      @              @      �?              $@      �?      @              @      �?              �?      @             @P@     �r@     �C@      q@      5@      j@      2@      j@      @      .@      @      @               @      @      �?              �?      @              @      (@      @      �?      @                      �?              &@      &@      h@      @      D@       @     �B@              6@       @      .@              "@       @      @      �?      @      �?      @      �?                      @              �?      �?              @      @      @                      @      @      c@      @     �@@              (@      @      5@      @      $@       @      $@       @       @              �?       @      �?              �?       @                       @       @                      &@      �?      ^@      �?      0@      �?      @              @      �?                      (@              Z@      @      �?              �?      @              2@     �O@      @     �I@      �?       @      �?                       @      @     �H@      �?       @               @      �?              @     �G@      �?      @              @      �?               @      F@      �?      C@              =@      �?      "@      �?       @               @      �?                      @      �?      @      �?       @      �?                       @              @      *@      (@      &@      @      �?      @              @      �?              $@      �?              �?      $@               @       @      �?              �?       @      �?       @      �?      �?              �?      �?                      �?              @      :@      >@              @      :@      8@      (@              ,@      8@      @      3@       @               @      3@      �?      �?              �?      �?              �?      2@              $@      �?       @              @      �?      �?      �?                      �?      $@      @      @      �?      @                      �?      @      @      �?      @              @      �?               @        �t�bub�       hhubehhub.